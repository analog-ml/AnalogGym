.param W_NM0=13 L_NM0=2 M_NM0=100
.param W_NM1=13 L_NM1=2 M_NM1=13
.param W_NM2=1 L_NM2=15 M_NM2=200
.param W_NM3=100 L_NM3=1 M_NM3=1
.param W_NM4=W_NM3 L_NM4=L_NM3 M_NM4=M_NM3
.param W_NM6=13 L_NM6=2 M_NM6=100
.param W_NM7=13 L_NM7=2 M_NM7=34
.param W_NM8=20 L_NM8=12 M_NM8=1
.param W_NM9=W_NM8 L_NM9=L_NM8 M_NM9=M_NM8
.param W_NM10=20 L_NM10=15 M_NM10=100
.param W_PM0=1.5 L_PM0=2 M_PM0=50
.param W_PM1=1.5 L_PM1=2 M_PM1=1
.param W_PM2=20 L_PM2=1 M_PM2=55
.param W_PM3=1.29 L_PM3=1.86 M_PM3=100
.param W_PM4=100 L_PM4=1 M_PM4=150
.param W_PM5=20 L_PM5=2 M_PM5=100
.param W_PM6=9 L_PM6=2 M_PM6=100
.param W_PM7=20 L_PM7=12 M_PM7=40
.param W_PM8=10 L_PM8=0.5 M_PM8=100
.param W_PM9=W_PM8 L_PM9=L_PM8 M_PM9=M_PM8
.param current_0_bias=5e-07
.param M_R0=100
.param M_C0=200
.param M_C1=160
.param M_C4=1
.param M_CL=5
