.param W_M0=3 L_M0=1 M_M0=1
.param W_M1=W_M0 L_M1=L_M0 M_M1=M_M0
.param W_M2=20 L_M2=4 M_M2=1
.param W_M3=W_M2 L_M3=L_M2 M_M3=M_M2
.param W_M4=1 L_M4=0.5 M_M4=1
.param W_M5=W_M4 L_M5=L_M4 M_M5=M_M4
.param W_M6=25 L_M6=1 M_M6=1
.param W_M7=3 L_M7=0.5 M_M7=1
.param W_M8=100 L_M8=1 M_M8=120
.param current_0_bias=5e-06
.param M_CL=200