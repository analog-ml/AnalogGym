let gmbs_NM0=@m.x1.XNM0.msky130_fd_pr__nfet_01v8[gmbs]
let gm_NM0=@m.x1.XNM0.msky130_fd_pr__nfet_01v8[gm]
let gds_NM0=@m.x1.XNM0.msky130_fd_pr__nfet_01v8[gds]
let vdsat_NM0=@m.x1.XNM0.msky130_fd_pr__nfet_01v8[vdsat]
let vth_NM0=@m.x1.XNM0.msky130_fd_pr__nfet_01v8[vth]
let id_NM0=@m.x1.XNM0.msky130_fd_pr__nfet_01v8[id]
let ibd_NM0=@m.x1.XNM0.msky130_fd_pr__nfet_01v8[ibd]
let ibs_NM0=@m.x1.XNM0.msky130_fd_pr__nfet_01v8[ibs]
let gbd_NM0=@m.x1.XNM0.msky130_fd_pr__nfet_01v8[gbd]
let gbs_NM0=@m.x1.XNM0.msky130_fd_pr__nfet_01v8[gbs]
let isub_NM0=@m.x1.XNM0.msky130_fd_pr__nfet_01v8[isub]
let igidl_NM0=@m.x1.XNM0.msky130_fd_pr__nfet_01v8[igidl]
let igisl_NM0=@m.x1.XNM0.msky130_fd_pr__nfet_01v8[igisl]
let igs_NM0=@m.x1.XNM0.msky130_fd_pr__nfet_01v8[igs]
let igd_NM0=@m.x1.XNM0.msky130_fd_pr__nfet_01v8[igd]
let igb_NM0=@m.x1.XNM0.msky130_fd_pr__nfet_01v8[igb]
let igcs_NM0=@m.x1.XNM0.msky130_fd_pr__nfet_01v8[igcs]
let vbs_NM0=@m.x1.XNM0.msky130_fd_pr__nfet_01v8[vbs]
let vgs_NM0=@m.x1.XNM0.msky130_fd_pr__nfet_01v8[vgs]
let vds_NM0=@m.x1.XNM0.msky130_fd_pr__nfet_01v8[vds]
let cgg_NM0=@m.x1.XNM0.msky130_fd_pr__nfet_01v8[cgg]
let cgs_NM0=@m.x1.XNM0.msky130_fd_pr__nfet_01v8[cgs]
let cgd_NM0=@m.x1.XNM0.msky130_fd_pr__nfet_01v8[cgd]
let cbg_NM0=@m.x1.XNM0.msky130_fd_pr__nfet_01v8[cbg]
let cbd_NM0=@m.x1.XNM0.msky130_fd_pr__nfet_01v8[cbd]
let cbs_NM0=@m.x1.XNM0.msky130_fd_pr__nfet_01v8[cbs]
let cdg_NM0=@m.x1.XNM0.msky130_fd_pr__nfet_01v8[cdg]
let cdd_NM0=@m.x1.XNM0.msky130_fd_pr__nfet_01v8[cdd]
let cds_NM0=@m.x1.XNM0.msky130_fd_pr__nfet_01v8[cds]
let csg_NM0=@m.x1.XNM0.msky130_fd_pr__nfet_01v8[csg]
let csd_NM0=@m.x1.XNM0.msky130_fd_pr__nfet_01v8[csd]
let css_NM0=@m.x1.XNM0.msky130_fd_pr__nfet_01v8[css]
let cgb_NM0=@m.x1.XNM0.msky130_fd_pr__nfet_01v8[cgb]
let cdb_NM0=@m.x1.XNM0.msky130_fd_pr__nfet_01v8[cdb]
let csb_NM0=@m.x1.XNM0.msky130_fd_pr__nfet_01v8[csb]
let cbb_NM0=@m.x1.XNM0.msky130_fd_pr__nfet_01v8[cbb]
let capbd_NM0=@m.x1.XNM0.msky130_fd_pr__nfet_01v8[capbd]
let capbs_NM0=@m.x1.XNM0.msky130_fd_pr__nfet_01v8[capbs]
let qg_NM0=@m.x1.XNM0.msky130_fd_pr__nfet_01v8[qg]
let qb_NM0=@m.x1.XNM0.msky130_fd_pr__nfet_01v8[qb]
let qs_NM0=@m.x1.XNM0.msky130_fd_pr__nfet_01v8[qs]
let qinv_NM0=@m.x1.XNM0.msky130_fd_pr__nfet_01v8[qinv]
let qdef_NM0=@m.x1.XNM0.msky130_fd_pr__nfet_01v8[qdef]
let gcrg_NM0=@m.x1.XNM0.msky130_fd_pr__nfet_01v8[gcrg]
let gtau_NM0=@m.x1.XNM0.msky130_fd_pr__nfet_01v8[gtau]

let gmbs_NM1=@m.x1.XNM1.msky130_fd_pr__nfet_01v8[gmbs]
let gm_NM1=@m.x1.XNM1.msky130_fd_pr__nfet_01v8[gm]
let gds_NM1=@m.x1.XNM1.msky130_fd_pr__nfet_01v8[gds]
let vdsat_NM1=@m.x1.XNM1.msky130_fd_pr__nfet_01v8[vdsat]
let vth_NM1=@m.x1.XNM1.msky130_fd_pr__nfet_01v8[vth]
let id_NM1=@m.x1.XNM1.msky130_fd_pr__nfet_01v8[id]
let ibd_NM1=@m.x1.XNM1.msky130_fd_pr__nfet_01v8[ibd]
let ibs_NM1=@m.x1.XNM1.msky130_fd_pr__nfet_01v8[ibs]
let gbd_NM1=@m.x1.XNM1.msky130_fd_pr__nfet_01v8[gbd]
let gbs_NM1=@m.x1.XNM1.msky130_fd_pr__nfet_01v8[gbs]
let isub_NM1=@m.x1.XNM1.msky130_fd_pr__nfet_01v8[isub]
let igidl_NM1=@m.x1.XNM1.msky130_fd_pr__nfet_01v8[igidl]
let igisl_NM1=@m.x1.XNM1.msky130_fd_pr__nfet_01v8[igisl]
let igs_NM1=@m.x1.XNM1.msky130_fd_pr__nfet_01v8[igs]
let igd_NM1=@m.x1.XNM1.msky130_fd_pr__nfet_01v8[igd]
let igb_NM1=@m.x1.XNM1.msky130_fd_pr__nfet_01v8[igb]
let igcs_NM1=@m.x1.XNM1.msky130_fd_pr__nfet_01v8[igcs]
let vbs_NM1=@m.x1.XNM1.msky130_fd_pr__nfet_01v8[vbs]
let vgs_NM1=@m.x1.XNM1.msky130_fd_pr__nfet_01v8[vgs]
let vds_NM1=@m.x1.XNM1.msky130_fd_pr__nfet_01v8[vds]
let cgg_NM1=@m.x1.XNM1.msky130_fd_pr__nfet_01v8[cgg]
let cgs_NM1=@m.x1.XNM1.msky130_fd_pr__nfet_01v8[cgs]
let cgd_NM1=@m.x1.XNM1.msky130_fd_pr__nfet_01v8[cgd]
let cbg_NM1=@m.x1.XNM1.msky130_fd_pr__nfet_01v8[cbg]
let cbd_NM1=@m.x1.XNM1.msky130_fd_pr__nfet_01v8[cbd]
let cbs_NM1=@m.x1.XNM1.msky130_fd_pr__nfet_01v8[cbs]
let cdg_NM1=@m.x1.XNM1.msky130_fd_pr__nfet_01v8[cdg]
let cdd_NM1=@m.x1.XNM1.msky130_fd_pr__nfet_01v8[cdd]
let cds_NM1=@m.x1.XNM1.msky130_fd_pr__nfet_01v8[cds]
let csg_NM1=@m.x1.XNM1.msky130_fd_pr__nfet_01v8[csg]
let csd_NM1=@m.x1.XNM1.msky130_fd_pr__nfet_01v8[csd]
let css_NM1=@m.x1.XNM1.msky130_fd_pr__nfet_01v8[css]
let cgb_NM1=@m.x1.XNM1.msky130_fd_pr__nfet_01v8[cgb]
let cdb_NM1=@m.x1.XNM1.msky130_fd_pr__nfet_01v8[cdb]
let csb_NM1=@m.x1.XNM1.msky130_fd_pr__nfet_01v8[csb]
let cbb_NM1=@m.x1.XNM1.msky130_fd_pr__nfet_01v8[cbb]
let capbd_NM1=@m.x1.XNM1.msky130_fd_pr__nfet_01v8[capbd]
let capbs_NM1=@m.x1.XNM1.msky130_fd_pr__nfet_01v8[capbs]
let qg_NM1=@m.x1.XNM1.msky130_fd_pr__nfet_01v8[qg]
let qb_NM1=@m.x1.XNM1.msky130_fd_pr__nfet_01v8[qb]
let qs_NM1=@m.x1.XNM1.msky130_fd_pr__nfet_01v8[qs]
let qinv_NM1=@m.x1.XNM1.msky130_fd_pr__nfet_01v8[qinv]
let qdef_NM1=@m.x1.XNM1.msky130_fd_pr__nfet_01v8[qdef]
let gcrg_NM1=@m.x1.XNM1.msky130_fd_pr__nfet_01v8[gcrg]
let gtau_NM1=@m.x1.XNM1.msky130_fd_pr__nfet_01v8[gtau]

let gmbs_NM2=@m.x1.XNM2.msky130_fd_pr__nfet_01v8[gmbs]
let gm_NM2=@m.x1.XNM2.msky130_fd_pr__nfet_01v8[gm]
let gds_NM2=@m.x1.XNM2.msky130_fd_pr__nfet_01v8[gds]
let vdsat_NM2=@m.x1.XNM2.msky130_fd_pr__nfet_01v8[vdsat]
let vth_NM2=@m.x1.XNM2.msky130_fd_pr__nfet_01v8[vth]
let id_NM2=@m.x1.XNM2.msky130_fd_pr__nfet_01v8[id]
let ibd_NM2=@m.x1.XNM2.msky130_fd_pr__nfet_01v8[ibd]
let ibs_NM2=@m.x1.XNM2.msky130_fd_pr__nfet_01v8[ibs]
let gbd_NM2=@m.x1.XNM2.msky130_fd_pr__nfet_01v8[gbd]
let gbs_NM2=@m.x1.XNM2.msky130_fd_pr__nfet_01v8[gbs]
let isub_NM2=@m.x1.XNM2.msky130_fd_pr__nfet_01v8[isub]
let igidl_NM2=@m.x1.XNM2.msky130_fd_pr__nfet_01v8[igidl]
let igisl_NM2=@m.x1.XNM2.msky130_fd_pr__nfet_01v8[igisl]
let igs_NM2=@m.x1.XNM2.msky130_fd_pr__nfet_01v8[igs]
let igd_NM2=@m.x1.XNM2.msky130_fd_pr__nfet_01v8[igd]
let igb_NM2=@m.x1.XNM2.msky130_fd_pr__nfet_01v8[igb]
let igcs_NM2=@m.x1.XNM2.msky130_fd_pr__nfet_01v8[igcs]
let vbs_NM2=@m.x1.XNM2.msky130_fd_pr__nfet_01v8[vbs]
let vgs_NM2=@m.x1.XNM2.msky130_fd_pr__nfet_01v8[vgs]
let vds_NM2=@m.x1.XNM2.msky130_fd_pr__nfet_01v8[vds]
let cgg_NM2=@m.x1.XNM2.msky130_fd_pr__nfet_01v8[cgg]
let cgs_NM2=@m.x1.XNM2.msky130_fd_pr__nfet_01v8[cgs]
let cgd_NM2=@m.x1.XNM2.msky130_fd_pr__nfet_01v8[cgd]
let cbg_NM2=@m.x1.XNM2.msky130_fd_pr__nfet_01v8[cbg]
let cbd_NM2=@m.x1.XNM2.msky130_fd_pr__nfet_01v8[cbd]
let cbs_NM2=@m.x1.XNM2.msky130_fd_pr__nfet_01v8[cbs]
let cdg_NM2=@m.x1.XNM2.msky130_fd_pr__nfet_01v8[cdg]
let cdd_NM2=@m.x1.XNM2.msky130_fd_pr__nfet_01v8[cdd]
let cds_NM2=@m.x1.XNM2.msky130_fd_pr__nfet_01v8[cds]
let csg_NM2=@m.x1.XNM2.msky130_fd_pr__nfet_01v8[csg]
let csd_NM2=@m.x1.XNM2.msky130_fd_pr__nfet_01v8[csd]
let css_NM2=@m.x1.XNM2.msky130_fd_pr__nfet_01v8[css]
let cgb_NM2=@m.x1.XNM2.msky130_fd_pr__nfet_01v8[cgb]
let cdb_NM2=@m.x1.XNM2.msky130_fd_pr__nfet_01v8[cdb]
let csb_NM2=@m.x1.XNM2.msky130_fd_pr__nfet_01v8[csb]
let cbb_NM2=@m.x1.XNM2.msky130_fd_pr__nfet_01v8[cbb]
let capbd_NM2=@m.x1.XNM2.msky130_fd_pr__nfet_01v8[capbd]
let capbs_NM2=@m.x1.XNM2.msky130_fd_pr__nfet_01v8[capbs]
let qg_NM2=@m.x1.XNM2.msky130_fd_pr__nfet_01v8[qg]
let qb_NM2=@m.x1.XNM2.msky130_fd_pr__nfet_01v8[qb]
let qs_NM2=@m.x1.XNM2.msky130_fd_pr__nfet_01v8[qs]
let qinv_NM2=@m.x1.XNM2.msky130_fd_pr__nfet_01v8[qinv]
let qdef_NM2=@m.x1.XNM2.msky130_fd_pr__nfet_01v8[qdef]
let gcrg_NM2=@m.x1.XNM2.msky130_fd_pr__nfet_01v8[gcrg]
let gtau_NM2=@m.x1.XNM2.msky130_fd_pr__nfet_01v8[gtau]

let gmbs_NM3=@m.x1.XNM3.msky130_fd_pr__nfet_01v8[gmbs]
let gm_NM3=@m.x1.XNM3.msky130_fd_pr__nfet_01v8[gm]
let gds_NM3=@m.x1.XNM3.msky130_fd_pr__nfet_01v8[gds]
let vdsat_NM3=@m.x1.XNM3.msky130_fd_pr__nfet_01v8[vdsat]
let vth_NM3=@m.x1.XNM3.msky130_fd_pr__nfet_01v8[vth]
let id_NM3=@m.x1.XNM3.msky130_fd_pr__nfet_01v8[id]
let ibd_NM3=@m.x1.XNM3.msky130_fd_pr__nfet_01v8[ibd]
let ibs_NM3=@m.x1.XNM3.msky130_fd_pr__nfet_01v8[ibs]
let gbd_NM3=@m.x1.XNM3.msky130_fd_pr__nfet_01v8[gbd]
let gbs_NM3=@m.x1.XNM3.msky130_fd_pr__nfet_01v8[gbs]
let isub_NM3=@m.x1.XNM3.msky130_fd_pr__nfet_01v8[isub]
let igidl_NM3=@m.x1.XNM3.msky130_fd_pr__nfet_01v8[igidl]
let igisl_NM3=@m.x1.XNM3.msky130_fd_pr__nfet_01v8[igisl]
let igs_NM3=@m.x1.XNM3.msky130_fd_pr__nfet_01v8[igs]
let igd_NM3=@m.x1.XNM3.msky130_fd_pr__nfet_01v8[igd]
let igb_NM3=@m.x1.XNM3.msky130_fd_pr__nfet_01v8[igb]
let igcs_NM3=@m.x1.XNM3.msky130_fd_pr__nfet_01v8[igcs]
let vbs_NM3=@m.x1.XNM3.msky130_fd_pr__nfet_01v8[vbs]
let vgs_NM3=@m.x1.XNM3.msky130_fd_pr__nfet_01v8[vgs]
let vds_NM3=@m.x1.XNM3.msky130_fd_pr__nfet_01v8[vds]
let cgg_NM3=@m.x1.XNM3.msky130_fd_pr__nfet_01v8[cgg]
let cgs_NM3=@m.x1.XNM3.msky130_fd_pr__nfet_01v8[cgs]
let cgd_NM3=@m.x1.XNM3.msky130_fd_pr__nfet_01v8[cgd]
let cbg_NM3=@m.x1.XNM3.msky130_fd_pr__nfet_01v8[cbg]
let cbd_NM3=@m.x1.XNM3.msky130_fd_pr__nfet_01v8[cbd]
let cbs_NM3=@m.x1.XNM3.msky130_fd_pr__nfet_01v8[cbs]
let cdg_NM3=@m.x1.XNM3.msky130_fd_pr__nfet_01v8[cdg]
let cdd_NM3=@m.x1.XNM3.msky130_fd_pr__nfet_01v8[cdd]
let cds_NM3=@m.x1.XNM3.msky130_fd_pr__nfet_01v8[cds]
let csg_NM3=@m.x1.XNM3.msky130_fd_pr__nfet_01v8[csg]
let csd_NM3=@m.x1.XNM3.msky130_fd_pr__nfet_01v8[csd]
let css_NM3=@m.x1.XNM3.msky130_fd_pr__nfet_01v8[css]
let cgb_NM3=@m.x1.XNM3.msky130_fd_pr__nfet_01v8[cgb]
let cdb_NM3=@m.x1.XNM3.msky130_fd_pr__nfet_01v8[cdb]
let csb_NM3=@m.x1.XNM3.msky130_fd_pr__nfet_01v8[csb]
let cbb_NM3=@m.x1.XNM3.msky130_fd_pr__nfet_01v8[cbb]
let capbd_NM3=@m.x1.XNM3.msky130_fd_pr__nfet_01v8[capbd]
let capbs_NM3=@m.x1.XNM3.msky130_fd_pr__nfet_01v8[capbs]
let qg_NM3=@m.x1.XNM3.msky130_fd_pr__nfet_01v8[qg]
let qb_NM3=@m.x1.XNM3.msky130_fd_pr__nfet_01v8[qb]
let qs_NM3=@m.x1.XNM3.msky130_fd_pr__nfet_01v8[qs]
let qinv_NM3=@m.x1.XNM3.msky130_fd_pr__nfet_01v8[qinv]
let qdef_NM3=@m.x1.XNM3.msky130_fd_pr__nfet_01v8[qdef]
let gcrg_NM3=@m.x1.XNM3.msky130_fd_pr__nfet_01v8[gcrg]
let gtau_NM3=@m.x1.XNM3.msky130_fd_pr__nfet_01v8[gtau]

let gmbs_NM4=@m.x1.XNM4.msky130_fd_pr__nfet_01v8[gmbs]
let gm_NM4=@m.x1.XNM4.msky130_fd_pr__nfet_01v8[gm]
let gds_NM4=@m.x1.XNM4.msky130_fd_pr__nfet_01v8[gds]
let vdsat_NM4=@m.x1.XNM4.msky130_fd_pr__nfet_01v8[vdsat]
let vth_NM4=@m.x1.XNM4.msky130_fd_pr__nfet_01v8[vth]
let id_NM4=@m.x1.XNM4.msky130_fd_pr__nfet_01v8[id]
let ibd_NM4=@m.x1.XNM4.msky130_fd_pr__nfet_01v8[ibd]
let ibs_NM4=@m.x1.XNM4.msky130_fd_pr__nfet_01v8[ibs]
let gbd_NM4=@m.x1.XNM4.msky130_fd_pr__nfet_01v8[gbd]
let gbs_NM4=@m.x1.XNM4.msky130_fd_pr__nfet_01v8[gbs]
let isub_NM4=@m.x1.XNM4.msky130_fd_pr__nfet_01v8[isub]
let igidl_NM4=@m.x1.XNM4.msky130_fd_pr__nfet_01v8[igidl]
let igisl_NM4=@m.x1.XNM4.msky130_fd_pr__nfet_01v8[igisl]
let igs_NM4=@m.x1.XNM4.msky130_fd_pr__nfet_01v8[igs]
let igd_NM4=@m.x1.XNM4.msky130_fd_pr__nfet_01v8[igd]
let igb_NM4=@m.x1.XNM4.msky130_fd_pr__nfet_01v8[igb]
let igcs_NM4=@m.x1.XNM4.msky130_fd_pr__nfet_01v8[igcs]
let vbs_NM4=@m.x1.XNM4.msky130_fd_pr__nfet_01v8[vbs]
let vgs_NM4=@m.x1.XNM4.msky130_fd_pr__nfet_01v8[vgs]
let vds_NM4=@m.x1.XNM4.msky130_fd_pr__nfet_01v8[vds]
let cgg_NM4=@m.x1.XNM4.msky130_fd_pr__nfet_01v8[cgg]
let cgs_NM4=@m.x1.XNM4.msky130_fd_pr__nfet_01v8[cgs]
let cgd_NM4=@m.x1.XNM4.msky130_fd_pr__nfet_01v8[cgd]
let cbg_NM4=@m.x1.XNM4.msky130_fd_pr__nfet_01v8[cbg]
let cbd_NM4=@m.x1.XNM4.msky130_fd_pr__nfet_01v8[cbd]
let cbs_NM4=@m.x1.XNM4.msky130_fd_pr__nfet_01v8[cbs]
let cdg_NM4=@m.x1.XNM4.msky130_fd_pr__nfet_01v8[cdg]
let cdd_NM4=@m.x1.XNM4.msky130_fd_pr__nfet_01v8[cdd]
let cds_NM4=@m.x1.XNM4.msky130_fd_pr__nfet_01v8[cds]
let csg_NM4=@m.x1.XNM4.msky130_fd_pr__nfet_01v8[csg]
let csd_NM4=@m.x1.XNM4.msky130_fd_pr__nfet_01v8[csd]
let css_NM4=@m.x1.XNM4.msky130_fd_pr__nfet_01v8[css]
let cgb_NM4=@m.x1.XNM4.msky130_fd_pr__nfet_01v8[cgb]
let cdb_NM4=@m.x1.XNM4.msky130_fd_pr__nfet_01v8[cdb]
let csb_NM4=@m.x1.XNM4.msky130_fd_pr__nfet_01v8[csb]
let cbb_NM4=@m.x1.XNM4.msky130_fd_pr__nfet_01v8[cbb]
let capbd_NM4=@m.x1.XNM4.msky130_fd_pr__nfet_01v8[capbd]
let capbs_NM4=@m.x1.XNM4.msky130_fd_pr__nfet_01v8[capbs]
let qg_NM4=@m.x1.XNM4.msky130_fd_pr__nfet_01v8[qg]
let qb_NM4=@m.x1.XNM4.msky130_fd_pr__nfet_01v8[qb]
let qs_NM4=@m.x1.XNM4.msky130_fd_pr__nfet_01v8[qs]
let qinv_NM4=@m.x1.XNM4.msky130_fd_pr__nfet_01v8[qinv]
let qdef_NM4=@m.x1.XNM4.msky130_fd_pr__nfet_01v8[qdef]
let gcrg_NM4=@m.x1.XNM4.msky130_fd_pr__nfet_01v8[gcrg]
let gtau_NM4=@m.x1.XNM4.msky130_fd_pr__nfet_01v8[gtau]

let gmbs_NM6=@m.x1.XNM6.msky130_fd_pr__nfet_01v8[gmbs]
let gm_NM6=@m.x1.XNM6.msky130_fd_pr__nfet_01v8[gm]
let gds_NM6=@m.x1.XNM6.msky130_fd_pr__nfet_01v8[gds]
let vdsat_NM6=@m.x1.XNM6.msky130_fd_pr__nfet_01v8[vdsat]
let vth_NM6=@m.x1.XNM6.msky130_fd_pr__nfet_01v8[vth]
let id_NM6=@m.x1.XNM6.msky130_fd_pr__nfet_01v8[id]
let ibd_NM6=@m.x1.XNM6.msky130_fd_pr__nfet_01v8[ibd]
let ibs_NM6=@m.x1.XNM6.msky130_fd_pr__nfet_01v8[ibs]
let gbd_NM6=@m.x1.XNM6.msky130_fd_pr__nfet_01v8[gbd]
let gbs_NM6=@m.x1.XNM6.msky130_fd_pr__nfet_01v8[gbs]
let isub_NM6=@m.x1.XNM6.msky130_fd_pr__nfet_01v8[isub]
let igidl_NM6=@m.x1.XNM6.msky130_fd_pr__nfet_01v8[igidl]
let igisl_NM6=@m.x1.XNM6.msky130_fd_pr__nfet_01v8[igisl]
let igs_NM6=@m.x1.XNM6.msky130_fd_pr__nfet_01v8[igs]
let igd_NM6=@m.x1.XNM6.msky130_fd_pr__nfet_01v8[igd]
let igb_NM6=@m.x1.XNM6.msky130_fd_pr__nfet_01v8[igb]
let igcs_NM6=@m.x1.XNM6.msky130_fd_pr__nfet_01v8[igcs]
let vbs_NM6=@m.x1.XNM6.msky130_fd_pr__nfet_01v8[vbs]
let vgs_NM6=@m.x1.XNM6.msky130_fd_pr__nfet_01v8[vgs]
let vds_NM6=@m.x1.XNM6.msky130_fd_pr__nfet_01v8[vds]
let cgg_NM6=@m.x1.XNM6.msky130_fd_pr__nfet_01v8[cgg]
let cgs_NM6=@m.x1.XNM6.msky130_fd_pr__nfet_01v8[cgs]
let cgd_NM6=@m.x1.XNM6.msky130_fd_pr__nfet_01v8[cgd]
let cbg_NM6=@m.x1.XNM6.msky130_fd_pr__nfet_01v8[cbg]
let cbd_NM6=@m.x1.XNM6.msky130_fd_pr__nfet_01v8[cbd]
let cbs_NM6=@m.x1.XNM6.msky130_fd_pr__nfet_01v8[cbs]
let cdg_NM6=@m.x1.XNM6.msky130_fd_pr__nfet_01v8[cdg]
let cdd_NM6=@m.x1.XNM6.msky130_fd_pr__nfet_01v8[cdd]
let cds_NM6=@m.x1.XNM6.msky130_fd_pr__nfet_01v8[cds]
let csg_NM6=@m.x1.XNM6.msky130_fd_pr__nfet_01v8[csg]
let csd_NM6=@m.x1.XNM6.msky130_fd_pr__nfet_01v8[csd]
let css_NM6=@m.x1.XNM6.msky130_fd_pr__nfet_01v8[css]
let cgb_NM6=@m.x1.XNM6.msky130_fd_pr__nfet_01v8[cgb]
let cdb_NM6=@m.x1.XNM6.msky130_fd_pr__nfet_01v8[cdb]
let csb_NM6=@m.x1.XNM6.msky130_fd_pr__nfet_01v8[csb]
let cbb_NM6=@m.x1.XNM6.msky130_fd_pr__nfet_01v8[cbb]
let capbd_NM6=@m.x1.XNM6.msky130_fd_pr__nfet_01v8[capbd]
let capbs_NM6=@m.x1.XNM6.msky130_fd_pr__nfet_01v8[capbs]
let qg_NM6=@m.x1.XNM6.msky130_fd_pr__nfet_01v8[qg]
let qb_NM6=@m.x1.XNM6.msky130_fd_pr__nfet_01v8[qb]
let qs_NM6=@m.x1.XNM6.msky130_fd_pr__nfet_01v8[qs]
let qinv_NM6=@m.x1.XNM6.msky130_fd_pr__nfet_01v8[qinv]
let qdef_NM6=@m.x1.XNM6.msky130_fd_pr__nfet_01v8[qdef]
let gcrg_NM6=@m.x1.XNM6.msky130_fd_pr__nfet_01v8[gcrg]
let gtau_NM6=@m.x1.XNM6.msky130_fd_pr__nfet_01v8[gtau]

let gmbs_NM7=@m.x1.XNM7.msky130_fd_pr__nfet_01v8[gmbs]
let gm_NM7=@m.x1.XNM7.msky130_fd_pr__nfet_01v8[gm]
let gds_NM7=@m.x1.XNM7.msky130_fd_pr__nfet_01v8[gds]
let vdsat_NM7=@m.x1.XNM7.msky130_fd_pr__nfet_01v8[vdsat]
let vth_NM7=@m.x1.XNM7.msky130_fd_pr__nfet_01v8[vth]
let id_NM7=@m.x1.XNM7.msky130_fd_pr__nfet_01v8[id]
let ibd_NM7=@m.x1.XNM7.msky130_fd_pr__nfet_01v8[ibd]
let ibs_NM7=@m.x1.XNM7.msky130_fd_pr__nfet_01v8[ibs]
let gbd_NM7=@m.x1.XNM7.msky130_fd_pr__nfet_01v8[gbd]
let gbs_NM7=@m.x1.XNM7.msky130_fd_pr__nfet_01v8[gbs]
let isub_NM7=@m.x1.XNM7.msky130_fd_pr__nfet_01v8[isub]
let igidl_NM7=@m.x1.XNM7.msky130_fd_pr__nfet_01v8[igidl]
let igisl_NM7=@m.x1.XNM7.msky130_fd_pr__nfet_01v8[igisl]
let igs_NM7=@m.x1.XNM7.msky130_fd_pr__nfet_01v8[igs]
let igd_NM7=@m.x1.XNM7.msky130_fd_pr__nfet_01v8[igd]
let igb_NM7=@m.x1.XNM7.msky130_fd_pr__nfet_01v8[igb]
let igcs_NM7=@m.x1.XNM7.msky130_fd_pr__nfet_01v8[igcs]
let vbs_NM7=@m.x1.XNM7.msky130_fd_pr__nfet_01v8[vbs]
let vgs_NM7=@m.x1.XNM7.msky130_fd_pr__nfet_01v8[vgs]
let vds_NM7=@m.x1.XNM7.msky130_fd_pr__nfet_01v8[vds]
let cgg_NM7=@m.x1.XNM7.msky130_fd_pr__nfet_01v8[cgg]
let cgs_NM7=@m.x1.XNM7.msky130_fd_pr__nfet_01v8[cgs]
let cgd_NM7=@m.x1.XNM7.msky130_fd_pr__nfet_01v8[cgd]
let cbg_NM7=@m.x1.XNM7.msky130_fd_pr__nfet_01v8[cbg]
let cbd_NM7=@m.x1.XNM7.msky130_fd_pr__nfet_01v8[cbd]
let cbs_NM7=@m.x1.XNM7.msky130_fd_pr__nfet_01v8[cbs]
let cdg_NM7=@m.x1.XNM7.msky130_fd_pr__nfet_01v8[cdg]
let cdd_NM7=@m.x1.XNM7.msky130_fd_pr__nfet_01v8[cdd]
let cds_NM7=@m.x1.XNM7.msky130_fd_pr__nfet_01v8[cds]
let csg_NM7=@m.x1.XNM7.msky130_fd_pr__nfet_01v8[csg]
let csd_NM7=@m.x1.XNM7.msky130_fd_pr__nfet_01v8[csd]
let css_NM7=@m.x1.XNM7.msky130_fd_pr__nfet_01v8[css]
let cgb_NM7=@m.x1.XNM7.msky130_fd_pr__nfet_01v8[cgb]
let cdb_NM7=@m.x1.XNM7.msky130_fd_pr__nfet_01v8[cdb]
let csb_NM7=@m.x1.XNM7.msky130_fd_pr__nfet_01v8[csb]
let cbb_NM7=@m.x1.XNM7.msky130_fd_pr__nfet_01v8[cbb]
let capbd_NM7=@m.x1.XNM7.msky130_fd_pr__nfet_01v8[capbd]
let capbs_NM7=@m.x1.XNM7.msky130_fd_pr__nfet_01v8[capbs]
let qg_NM7=@m.x1.XNM7.msky130_fd_pr__nfet_01v8[qg]
let qb_NM7=@m.x1.XNM7.msky130_fd_pr__nfet_01v8[qb]
let qs_NM7=@m.x1.XNM7.msky130_fd_pr__nfet_01v8[qs]
let qinv_NM7=@m.x1.XNM7.msky130_fd_pr__nfet_01v8[qinv]
let qdef_NM7=@m.x1.XNM7.msky130_fd_pr__nfet_01v8[qdef]
let gcrg_NM7=@m.x1.XNM7.msky130_fd_pr__nfet_01v8[gcrg]
let gtau_NM7=@m.x1.XNM7.msky130_fd_pr__nfet_01v8[gtau]

let gmbs_NM8=@m.x1.XNM8.msky130_fd_pr__nfet_01v8[gmbs]
let gm_NM8=@m.x1.XNM8.msky130_fd_pr__nfet_01v8[gm]
let gds_NM8=@m.x1.XNM8.msky130_fd_pr__nfet_01v8[gds]
let vdsat_NM8=@m.x1.XNM8.msky130_fd_pr__nfet_01v8[vdsat]
let vth_NM8=@m.x1.XNM8.msky130_fd_pr__nfet_01v8[vth]
let id_NM8=@m.x1.XNM8.msky130_fd_pr__nfet_01v8[id]
let ibd_NM8=@m.x1.XNM8.msky130_fd_pr__nfet_01v8[ibd]
let ibs_NM8=@m.x1.XNM8.msky130_fd_pr__nfet_01v8[ibs]
let gbd_NM8=@m.x1.XNM8.msky130_fd_pr__nfet_01v8[gbd]
let gbs_NM8=@m.x1.XNM8.msky130_fd_pr__nfet_01v8[gbs]
let isub_NM8=@m.x1.XNM8.msky130_fd_pr__nfet_01v8[isub]
let igidl_NM8=@m.x1.XNM8.msky130_fd_pr__nfet_01v8[igidl]
let igisl_NM8=@m.x1.XNM8.msky130_fd_pr__nfet_01v8[igisl]
let igs_NM8=@m.x1.XNM8.msky130_fd_pr__nfet_01v8[igs]
let igd_NM8=@m.x1.XNM8.msky130_fd_pr__nfet_01v8[igd]
let igb_NM8=@m.x1.XNM8.msky130_fd_pr__nfet_01v8[igb]
let igcs_NM8=@m.x1.XNM8.msky130_fd_pr__nfet_01v8[igcs]
let vbs_NM8=@m.x1.XNM8.msky130_fd_pr__nfet_01v8[vbs]
let vgs_NM8=@m.x1.XNM8.msky130_fd_pr__nfet_01v8[vgs]
let vds_NM8=@m.x1.XNM8.msky130_fd_pr__nfet_01v8[vds]
let cgg_NM8=@m.x1.XNM8.msky130_fd_pr__nfet_01v8[cgg]
let cgs_NM8=@m.x1.XNM8.msky130_fd_pr__nfet_01v8[cgs]
let cgd_NM8=@m.x1.XNM8.msky130_fd_pr__nfet_01v8[cgd]
let cbg_NM8=@m.x1.XNM8.msky130_fd_pr__nfet_01v8[cbg]
let cbd_NM8=@m.x1.XNM8.msky130_fd_pr__nfet_01v8[cbd]
let cbs_NM8=@m.x1.XNM8.msky130_fd_pr__nfet_01v8[cbs]
let cdg_NM8=@m.x1.XNM8.msky130_fd_pr__nfet_01v8[cdg]
let cdd_NM8=@m.x1.XNM8.msky130_fd_pr__nfet_01v8[cdd]
let cds_NM8=@m.x1.XNM8.msky130_fd_pr__nfet_01v8[cds]
let csg_NM8=@m.x1.XNM8.msky130_fd_pr__nfet_01v8[csg]
let csd_NM8=@m.x1.XNM8.msky130_fd_pr__nfet_01v8[csd]
let css_NM8=@m.x1.XNM8.msky130_fd_pr__nfet_01v8[css]
let cgb_NM8=@m.x1.XNM8.msky130_fd_pr__nfet_01v8[cgb]
let cdb_NM8=@m.x1.XNM8.msky130_fd_pr__nfet_01v8[cdb]
let csb_NM8=@m.x1.XNM8.msky130_fd_pr__nfet_01v8[csb]
let cbb_NM8=@m.x1.XNM8.msky130_fd_pr__nfet_01v8[cbb]
let capbd_NM8=@m.x1.XNM8.msky130_fd_pr__nfet_01v8[capbd]
let capbs_NM8=@m.x1.XNM8.msky130_fd_pr__nfet_01v8[capbs]
let qg_NM8=@m.x1.XNM8.msky130_fd_pr__nfet_01v8[qg]
let qb_NM8=@m.x1.XNM8.msky130_fd_pr__nfet_01v8[qb]
let qs_NM8=@m.x1.XNM8.msky130_fd_pr__nfet_01v8[qs]
let qinv_NM8=@m.x1.XNM8.msky130_fd_pr__nfet_01v8[qinv]
let qdef_NM8=@m.x1.XNM8.msky130_fd_pr__nfet_01v8[qdef]
let gcrg_NM8=@m.x1.XNM8.msky130_fd_pr__nfet_01v8[gcrg]
let gtau_NM8=@m.x1.XNM8.msky130_fd_pr__nfet_01v8[gtau]

let gmbs_NM9=@m.x1.XNM9.msky130_fd_pr__nfet_01v8[gmbs]
let gm_NM9=@m.x1.XNM9.msky130_fd_pr__nfet_01v8[gm]
let gds_NM9=@m.x1.XNM9.msky130_fd_pr__nfet_01v8[gds]
let vdsat_NM9=@m.x1.XNM9.msky130_fd_pr__nfet_01v8[vdsat]
let vth_NM9=@m.x1.XNM9.msky130_fd_pr__nfet_01v8[vth]
let id_NM9=@m.x1.XNM9.msky130_fd_pr__nfet_01v8[id]
let ibd_NM9=@m.x1.XNM9.msky130_fd_pr__nfet_01v8[ibd]
let ibs_NM9=@m.x1.XNM9.msky130_fd_pr__nfet_01v8[ibs]
let gbd_NM9=@m.x1.XNM9.msky130_fd_pr__nfet_01v8[gbd]
let gbs_NM9=@m.x1.XNM9.msky130_fd_pr__nfet_01v8[gbs]
let isub_NM9=@m.x1.XNM9.msky130_fd_pr__nfet_01v8[isub]
let igidl_NM9=@m.x1.XNM9.msky130_fd_pr__nfet_01v8[igidl]
let igisl_NM9=@m.x1.XNM9.msky130_fd_pr__nfet_01v8[igisl]
let igs_NM9=@m.x1.XNM9.msky130_fd_pr__nfet_01v8[igs]
let igd_NM9=@m.x1.XNM9.msky130_fd_pr__nfet_01v8[igd]
let igb_NM9=@m.x1.XNM9.msky130_fd_pr__nfet_01v8[igb]
let igcs_NM9=@m.x1.XNM9.msky130_fd_pr__nfet_01v8[igcs]
let vbs_NM9=@m.x1.XNM9.msky130_fd_pr__nfet_01v8[vbs]
let vgs_NM9=@m.x1.XNM9.msky130_fd_pr__nfet_01v8[vgs]
let vds_NM9=@m.x1.XNM9.msky130_fd_pr__nfet_01v8[vds]
let cgg_NM9=@m.x1.XNM9.msky130_fd_pr__nfet_01v8[cgg]
let cgs_NM9=@m.x1.XNM9.msky130_fd_pr__nfet_01v8[cgs]
let cgd_NM9=@m.x1.XNM9.msky130_fd_pr__nfet_01v8[cgd]
let cbg_NM9=@m.x1.XNM9.msky130_fd_pr__nfet_01v8[cbg]
let cbd_NM9=@m.x1.XNM9.msky130_fd_pr__nfet_01v8[cbd]
let cbs_NM9=@m.x1.XNM9.msky130_fd_pr__nfet_01v8[cbs]
let cdg_NM9=@m.x1.XNM9.msky130_fd_pr__nfet_01v8[cdg]
let cdd_NM9=@m.x1.XNM9.msky130_fd_pr__nfet_01v8[cdd]
let cds_NM9=@m.x1.XNM9.msky130_fd_pr__nfet_01v8[cds]
let csg_NM9=@m.x1.XNM9.msky130_fd_pr__nfet_01v8[csg]
let csd_NM9=@m.x1.XNM9.msky130_fd_pr__nfet_01v8[csd]
let css_NM9=@m.x1.XNM9.msky130_fd_pr__nfet_01v8[css]
let cgb_NM9=@m.x1.XNM9.msky130_fd_pr__nfet_01v8[cgb]
let cdb_NM9=@m.x1.XNM9.msky130_fd_pr__nfet_01v8[cdb]
let csb_NM9=@m.x1.XNM9.msky130_fd_pr__nfet_01v8[csb]
let cbb_NM9=@m.x1.XNM9.msky130_fd_pr__nfet_01v8[cbb]
let capbd_NM9=@m.x1.XNM9.msky130_fd_pr__nfet_01v8[capbd]
let capbs_NM9=@m.x1.XNM9.msky130_fd_pr__nfet_01v8[capbs]
let qg_NM9=@m.x1.XNM9.msky130_fd_pr__nfet_01v8[qg]
let qb_NM9=@m.x1.XNM9.msky130_fd_pr__nfet_01v8[qb]
let qs_NM9=@m.x1.XNM9.msky130_fd_pr__nfet_01v8[qs]
let qinv_NM9=@m.x1.XNM9.msky130_fd_pr__nfet_01v8[qinv]
let qdef_NM9=@m.x1.XNM9.msky130_fd_pr__nfet_01v8[qdef]
let gcrg_NM9=@m.x1.XNM9.msky130_fd_pr__nfet_01v8[gcrg]
let gtau_NM9=@m.x1.XNM9.msky130_fd_pr__nfet_01v8[gtau]

let gmbs_NM10=@m.x1.XNM10.msky130_fd_pr__nfet_01v8[gmbs]
let gm_NM10=@m.x1.XNM10.msky130_fd_pr__nfet_01v8[gm]
let gds_NM10=@m.x1.XNM10.msky130_fd_pr__nfet_01v8[gds]
let vdsat_NM10=@m.x1.XNM10.msky130_fd_pr__nfet_01v8[vdsat]
let vth_NM10=@m.x1.XNM10.msky130_fd_pr__nfet_01v8[vth]
let id_NM10=@m.x1.XNM10.msky130_fd_pr__nfet_01v8[id]
let ibd_NM10=@m.x1.XNM10.msky130_fd_pr__nfet_01v8[ibd]
let ibs_NM10=@m.x1.XNM10.msky130_fd_pr__nfet_01v8[ibs]
let gbd_NM10=@m.x1.XNM10.msky130_fd_pr__nfet_01v8[gbd]
let gbs_NM10=@m.x1.XNM10.msky130_fd_pr__nfet_01v8[gbs]
let isub_NM10=@m.x1.XNM10.msky130_fd_pr__nfet_01v8[isub]
let igidl_NM10=@m.x1.XNM10.msky130_fd_pr__nfet_01v8[igidl]
let igisl_NM10=@m.x1.XNM10.msky130_fd_pr__nfet_01v8[igisl]
let igs_NM10=@m.x1.XNM10.msky130_fd_pr__nfet_01v8[igs]
let igd_NM10=@m.x1.XNM10.msky130_fd_pr__nfet_01v8[igd]
let igb_NM10=@m.x1.XNM10.msky130_fd_pr__nfet_01v8[igb]
let igcs_NM10=@m.x1.XNM10.msky130_fd_pr__nfet_01v8[igcs]
let vbs_NM10=@m.x1.XNM10.msky130_fd_pr__nfet_01v8[vbs]
let vgs_NM10=@m.x1.XNM10.msky130_fd_pr__nfet_01v8[vgs]
let vds_NM10=@m.x1.XNM10.msky130_fd_pr__nfet_01v8[vds]
let cgg_NM10=@m.x1.XNM10.msky130_fd_pr__nfet_01v8[cgg]
let cgs_NM10=@m.x1.XNM10.msky130_fd_pr__nfet_01v8[cgs]
let cgd_NM10=@m.x1.XNM10.msky130_fd_pr__nfet_01v8[cgd]
let cbg_NM10=@m.x1.XNM10.msky130_fd_pr__nfet_01v8[cbg]
let cbd_NM10=@m.x1.XNM10.msky130_fd_pr__nfet_01v8[cbd]
let cbs_NM10=@m.x1.XNM10.msky130_fd_pr__nfet_01v8[cbs]
let cdg_NM10=@m.x1.XNM10.msky130_fd_pr__nfet_01v8[cdg]
let cdd_NM10=@m.x1.XNM10.msky130_fd_pr__nfet_01v8[cdd]
let cds_NM10=@m.x1.XNM10.msky130_fd_pr__nfet_01v8[cds]
let csg_NM10=@m.x1.XNM10.msky130_fd_pr__nfet_01v8[csg]
let csd_NM10=@m.x1.XNM10.msky130_fd_pr__nfet_01v8[csd]
let css_NM10=@m.x1.XNM10.msky130_fd_pr__nfet_01v8[css]
let cgb_NM10=@m.x1.XNM10.msky130_fd_pr__nfet_01v8[cgb]
let cdb_NM10=@m.x1.XNM10.msky130_fd_pr__nfet_01v8[cdb]
let csb_NM10=@m.x1.XNM10.msky130_fd_pr__nfet_01v8[csb]
let cbb_NM10=@m.x1.XNM10.msky130_fd_pr__nfet_01v8[cbb]
let capbd_NM10=@m.x1.XNM10.msky130_fd_pr__nfet_01v8[capbd]
let capbs_NM10=@m.x1.XNM10.msky130_fd_pr__nfet_01v8[capbs]
let qg_NM10=@m.x1.XNM10.msky130_fd_pr__nfet_01v8[qg]
let qb_NM10=@m.x1.XNM10.msky130_fd_pr__nfet_01v8[qb]
let qs_NM10=@m.x1.XNM10.msky130_fd_pr__nfet_01v8[qs]
let qinv_NM10=@m.x1.XNM10.msky130_fd_pr__nfet_01v8[qinv]
let qdef_NM10=@m.x1.XNM10.msky130_fd_pr__nfet_01v8[qdef]
let gcrg_NM10=@m.x1.XNM10.msky130_fd_pr__nfet_01v8[gcrg]
let gtau_NM10=@m.x1.XNM10.msky130_fd_pr__nfet_01v8[gtau]

let gmbs_PM0=@m.x1.XPM0.msky130_fd_pr__pfet_01v8[gmbs]
let gm_PM0=@m.x1.XPM0.msky130_fd_pr__pfet_01v8[gm]
let gds_PM0=@m.x1.XPM0.msky130_fd_pr__pfet_01v8[gds]
let vdsat_PM0=@m.x1.XPM0.msky130_fd_pr__pfet_01v8[vdsat]
let vth_PM0=@m.x1.XPM0.msky130_fd_pr__pfet_01v8[vth]
let id_PM0=@m.x1.XPM0.msky130_fd_pr__pfet_01v8[id]
let ibd_PM0=@m.x1.XPM0.msky130_fd_pr__pfet_01v8[ibd]
let ibs_PM0=@m.x1.XPM0.msky130_fd_pr__pfet_01v8[ibs]
let gbd_PM0=@m.x1.XPM0.msky130_fd_pr__pfet_01v8[gbd]
let gbs_PM0=@m.x1.XPM0.msky130_fd_pr__pfet_01v8[gbs]
let isub_PM0=@m.x1.XPM0.msky130_fd_pr__pfet_01v8[isub]
let igidl_PM0=@m.x1.XPM0.msky130_fd_pr__pfet_01v8[igidl]
let igisl_PM0=@m.x1.XPM0.msky130_fd_pr__pfet_01v8[igisl]
let igs_PM0=@m.x1.XPM0.msky130_fd_pr__pfet_01v8[igs]
let igd_PM0=@m.x1.XPM0.msky130_fd_pr__pfet_01v8[igd]
let igb_PM0=@m.x1.XPM0.msky130_fd_pr__pfet_01v8[igb]
let igcs_PM0=@m.x1.XPM0.msky130_fd_pr__pfet_01v8[igcs]
let vbs_PM0=@m.x1.XPM0.msky130_fd_pr__pfet_01v8[vbs]
let vgs_PM0=@m.x1.XPM0.msky130_fd_pr__pfet_01v8[vgs]
let vds_PM0=@m.x1.XPM0.msky130_fd_pr__pfet_01v8[vds]
let cgg_PM0=@m.x1.XPM0.msky130_fd_pr__pfet_01v8[cgg]
let cgs_PM0=@m.x1.XPM0.msky130_fd_pr__pfet_01v8[cgs]
let cgd_PM0=@m.x1.XPM0.msky130_fd_pr__pfet_01v8[cgd]
let cbg_PM0=@m.x1.XPM0.msky130_fd_pr__pfet_01v8[cbg]
let cbd_PM0=@m.x1.XPM0.msky130_fd_pr__pfet_01v8[cbd]
let cbs_PM0=@m.x1.XPM0.msky130_fd_pr__pfet_01v8[cbs]
let cdg_PM0=@m.x1.XPM0.msky130_fd_pr__pfet_01v8[cdg]
let cdd_PM0=@m.x1.XPM0.msky130_fd_pr__pfet_01v8[cdd]
let cds_PM0=@m.x1.XPM0.msky130_fd_pr__pfet_01v8[cds]
let csg_PM0=@m.x1.XPM0.msky130_fd_pr__pfet_01v8[csg]
let csd_PM0=@m.x1.XPM0.msky130_fd_pr__pfet_01v8[csd]
let css_PM0=@m.x1.XPM0.msky130_fd_pr__pfet_01v8[css]
let cgb_PM0=@m.x1.XPM0.msky130_fd_pr__pfet_01v8[cgb]
let cdb_PM0=@m.x1.XPM0.msky130_fd_pr__pfet_01v8[cdb]
let csb_PM0=@m.x1.XPM0.msky130_fd_pr__pfet_01v8[csb]
let cbb_PM0=@m.x1.XPM0.msky130_fd_pr__pfet_01v8[cbb]
let capbd_PM0=@m.x1.XPM0.msky130_fd_pr__pfet_01v8[capbd]
let capbs_PM0=@m.x1.XPM0.msky130_fd_pr__pfet_01v8[capbs]
let qg_PM0=@m.x1.XPM0.msky130_fd_pr__pfet_01v8[qg]
let qb_PM0=@m.x1.XPM0.msky130_fd_pr__pfet_01v8[qb]
let qs_PM0=@m.x1.XPM0.msky130_fd_pr__pfet_01v8[qs]
let qinv_PM0=@m.x1.XPM0.msky130_fd_pr__pfet_01v8[qinv]
let qdef_PM0=@m.x1.XPM0.msky130_fd_pr__pfet_01v8[qdef]
let gcrg_PM0=@m.x1.XPM0.msky130_fd_pr__pfet_01v8[gcrg]
let gtau_PM0=@m.x1.XPM0.msky130_fd_pr__pfet_01v8[gtau]

let gmbs_PM1=@m.x1.XPM1.msky130_fd_pr__pfet_01v8[gmbs]
let gm_PM1=@m.x1.XPM1.msky130_fd_pr__pfet_01v8[gm]
let gds_PM1=@m.x1.XPM1.msky130_fd_pr__pfet_01v8[gds]
let vdsat_PM1=@m.x1.XPM1.msky130_fd_pr__pfet_01v8[vdsat]
let vth_PM1=@m.x1.XPM1.msky130_fd_pr__pfet_01v8[vth]
let id_PM1=@m.x1.XPM1.msky130_fd_pr__pfet_01v8[id]
let ibd_PM1=@m.x1.XPM1.msky130_fd_pr__pfet_01v8[ibd]
let ibs_PM1=@m.x1.XPM1.msky130_fd_pr__pfet_01v8[ibs]
let gbd_PM1=@m.x1.XPM1.msky130_fd_pr__pfet_01v8[gbd]
let gbs_PM1=@m.x1.XPM1.msky130_fd_pr__pfet_01v8[gbs]
let isub_PM1=@m.x1.XPM1.msky130_fd_pr__pfet_01v8[isub]
let igidl_PM1=@m.x1.XPM1.msky130_fd_pr__pfet_01v8[igidl]
let igisl_PM1=@m.x1.XPM1.msky130_fd_pr__pfet_01v8[igisl]
let igs_PM1=@m.x1.XPM1.msky130_fd_pr__pfet_01v8[igs]
let igd_PM1=@m.x1.XPM1.msky130_fd_pr__pfet_01v8[igd]
let igb_PM1=@m.x1.XPM1.msky130_fd_pr__pfet_01v8[igb]
let igcs_PM1=@m.x1.XPM1.msky130_fd_pr__pfet_01v8[igcs]
let vbs_PM1=@m.x1.XPM1.msky130_fd_pr__pfet_01v8[vbs]
let vgs_PM1=@m.x1.XPM1.msky130_fd_pr__pfet_01v8[vgs]
let vds_PM1=@m.x1.XPM1.msky130_fd_pr__pfet_01v8[vds]
let cgg_PM1=@m.x1.XPM1.msky130_fd_pr__pfet_01v8[cgg]
let cgs_PM1=@m.x1.XPM1.msky130_fd_pr__pfet_01v8[cgs]
let cgd_PM1=@m.x1.XPM1.msky130_fd_pr__pfet_01v8[cgd]
let cbg_PM1=@m.x1.XPM1.msky130_fd_pr__pfet_01v8[cbg]
let cbd_PM1=@m.x1.XPM1.msky130_fd_pr__pfet_01v8[cbd]
let cbs_PM1=@m.x1.XPM1.msky130_fd_pr__pfet_01v8[cbs]
let cdg_PM1=@m.x1.XPM1.msky130_fd_pr__pfet_01v8[cdg]
let cdd_PM1=@m.x1.XPM1.msky130_fd_pr__pfet_01v8[cdd]
let cds_PM1=@m.x1.XPM1.msky130_fd_pr__pfet_01v8[cds]
let csg_PM1=@m.x1.XPM1.msky130_fd_pr__pfet_01v8[csg]
let csd_PM1=@m.x1.XPM1.msky130_fd_pr__pfet_01v8[csd]
let css_PM1=@m.x1.XPM1.msky130_fd_pr__pfet_01v8[css]
let cgb_PM1=@m.x1.XPM1.msky130_fd_pr__pfet_01v8[cgb]
let cdb_PM1=@m.x1.XPM1.msky130_fd_pr__pfet_01v8[cdb]
let csb_PM1=@m.x1.XPM1.msky130_fd_pr__pfet_01v8[csb]
let cbb_PM1=@m.x1.XPM1.msky130_fd_pr__pfet_01v8[cbb]
let capbd_PM1=@m.x1.XPM1.msky130_fd_pr__pfet_01v8[capbd]
let capbs_PM1=@m.x1.XPM1.msky130_fd_pr__pfet_01v8[capbs]
let qg_PM1=@m.x1.XPM1.msky130_fd_pr__pfet_01v8[qg]
let qb_PM1=@m.x1.XPM1.msky130_fd_pr__pfet_01v8[qb]
let qs_PM1=@m.x1.XPM1.msky130_fd_pr__pfet_01v8[qs]
let qinv_PM1=@m.x1.XPM1.msky130_fd_pr__pfet_01v8[qinv]
let qdef_PM1=@m.x1.XPM1.msky130_fd_pr__pfet_01v8[qdef]
let gcrg_PM1=@m.x1.XPM1.msky130_fd_pr__pfet_01v8[gcrg]
let gtau_PM1=@m.x1.XPM1.msky130_fd_pr__pfet_01v8[gtau]

let gmbs_PM2=@m.x1.XPM2.msky130_fd_pr__pfet_01v8[gmbs]
let gm_PM2=@m.x1.XPM2.msky130_fd_pr__pfet_01v8[gm]
let gds_PM2=@m.x1.XPM2.msky130_fd_pr__pfet_01v8[gds]
let vdsat_PM2=@m.x1.XPM2.msky130_fd_pr__pfet_01v8[vdsat]
let vth_PM2=@m.x1.XPM2.msky130_fd_pr__pfet_01v8[vth]
let id_PM2=@m.x1.XPM2.msky130_fd_pr__pfet_01v8[id]
let ibd_PM2=@m.x1.XPM2.msky130_fd_pr__pfet_01v8[ibd]
let ibs_PM2=@m.x1.XPM2.msky130_fd_pr__pfet_01v8[ibs]
let gbd_PM2=@m.x1.XPM2.msky130_fd_pr__pfet_01v8[gbd]
let gbs_PM2=@m.x1.XPM2.msky130_fd_pr__pfet_01v8[gbs]
let isub_PM2=@m.x1.XPM2.msky130_fd_pr__pfet_01v8[isub]
let igidl_PM2=@m.x1.XPM2.msky130_fd_pr__pfet_01v8[igidl]
let igisl_PM2=@m.x1.XPM2.msky130_fd_pr__pfet_01v8[igisl]
let igs_PM2=@m.x1.XPM2.msky130_fd_pr__pfet_01v8[igs]
let igd_PM2=@m.x1.XPM2.msky130_fd_pr__pfet_01v8[igd]
let igb_PM2=@m.x1.XPM2.msky130_fd_pr__pfet_01v8[igb]
let igcs_PM2=@m.x1.XPM2.msky130_fd_pr__pfet_01v8[igcs]
let vbs_PM2=@m.x1.XPM2.msky130_fd_pr__pfet_01v8[vbs]
let vgs_PM2=@m.x1.XPM2.msky130_fd_pr__pfet_01v8[vgs]
let vds_PM2=@m.x1.XPM2.msky130_fd_pr__pfet_01v8[vds]
let cgg_PM2=@m.x1.XPM2.msky130_fd_pr__pfet_01v8[cgg]
let cgs_PM2=@m.x1.XPM2.msky130_fd_pr__pfet_01v8[cgs]
let cgd_PM2=@m.x1.XPM2.msky130_fd_pr__pfet_01v8[cgd]
let cbg_PM2=@m.x1.XPM2.msky130_fd_pr__pfet_01v8[cbg]
let cbd_PM2=@m.x1.XPM2.msky130_fd_pr__pfet_01v8[cbd]
let cbs_PM2=@m.x1.XPM2.msky130_fd_pr__pfet_01v8[cbs]
let cdg_PM2=@m.x1.XPM2.msky130_fd_pr__pfet_01v8[cdg]
let cdd_PM2=@m.x1.XPM2.msky130_fd_pr__pfet_01v8[cdd]
let cds_PM2=@m.x1.XPM2.msky130_fd_pr__pfet_01v8[cds]
let csg_PM2=@m.x1.XPM2.msky130_fd_pr__pfet_01v8[csg]
let csd_PM2=@m.x1.XPM2.msky130_fd_pr__pfet_01v8[csd]
let css_PM2=@m.x1.XPM2.msky130_fd_pr__pfet_01v8[css]
let cgb_PM2=@m.x1.XPM2.msky130_fd_pr__pfet_01v8[cgb]
let cdb_PM2=@m.x1.XPM2.msky130_fd_pr__pfet_01v8[cdb]
let csb_PM2=@m.x1.XPM2.msky130_fd_pr__pfet_01v8[csb]
let cbb_PM2=@m.x1.XPM2.msky130_fd_pr__pfet_01v8[cbb]
let capbd_PM2=@m.x1.XPM2.msky130_fd_pr__pfet_01v8[capbd]
let capbs_PM2=@m.x1.XPM2.msky130_fd_pr__pfet_01v8[capbs]
let qg_PM2=@m.x1.XPM2.msky130_fd_pr__pfet_01v8[qg]
let qb_PM2=@m.x1.XPM2.msky130_fd_pr__pfet_01v8[qb]
let qs_PM2=@m.x1.XPM2.msky130_fd_pr__pfet_01v8[qs]
let qinv_PM2=@m.x1.XPM2.msky130_fd_pr__pfet_01v8[qinv]
let qdef_PM2=@m.x1.XPM2.msky130_fd_pr__pfet_01v8[qdef]
let gcrg_PM2=@m.x1.XPM2.msky130_fd_pr__pfet_01v8[gcrg]
let gtau_PM2=@m.x1.XPM2.msky130_fd_pr__pfet_01v8[gtau]

let gmbs_PM3=@m.x1.XPM3.msky130_fd_pr__pfet_01v8[gmbs]
let gm_PM3=@m.x1.XPM3.msky130_fd_pr__pfet_01v8[gm]
let gds_PM3=@m.x1.XPM3.msky130_fd_pr__pfet_01v8[gds]
let vdsat_PM3=@m.x1.XPM3.msky130_fd_pr__pfet_01v8[vdsat]
let vth_PM3=@m.x1.XPM3.msky130_fd_pr__pfet_01v8[vth]
let id_PM3=@m.x1.XPM3.msky130_fd_pr__pfet_01v8[id]
let ibd_PM3=@m.x1.XPM3.msky130_fd_pr__pfet_01v8[ibd]
let ibs_PM3=@m.x1.XPM3.msky130_fd_pr__pfet_01v8[ibs]
let gbd_PM3=@m.x1.XPM3.msky130_fd_pr__pfet_01v8[gbd]
let gbs_PM3=@m.x1.XPM3.msky130_fd_pr__pfet_01v8[gbs]
let isub_PM3=@m.x1.XPM3.msky130_fd_pr__pfet_01v8[isub]
let igidl_PM3=@m.x1.XPM3.msky130_fd_pr__pfet_01v8[igidl]
let igisl_PM3=@m.x1.XPM3.msky130_fd_pr__pfet_01v8[igisl]
let igs_PM3=@m.x1.XPM3.msky130_fd_pr__pfet_01v8[igs]
let igd_PM3=@m.x1.XPM3.msky130_fd_pr__pfet_01v8[igd]
let igb_PM3=@m.x1.XPM3.msky130_fd_pr__pfet_01v8[igb]
let igcs_PM3=@m.x1.XPM3.msky130_fd_pr__pfet_01v8[igcs]
let vbs_PM3=@m.x1.XPM3.msky130_fd_pr__pfet_01v8[vbs]
let vgs_PM3=@m.x1.XPM3.msky130_fd_pr__pfet_01v8[vgs]
let vds_PM3=@m.x1.XPM3.msky130_fd_pr__pfet_01v8[vds]
let cgg_PM3=@m.x1.XPM3.msky130_fd_pr__pfet_01v8[cgg]
let cgs_PM3=@m.x1.XPM3.msky130_fd_pr__pfet_01v8[cgs]
let cgd_PM3=@m.x1.XPM3.msky130_fd_pr__pfet_01v8[cgd]
let cbg_PM3=@m.x1.XPM3.msky130_fd_pr__pfet_01v8[cbg]
let cbd_PM3=@m.x1.XPM3.msky130_fd_pr__pfet_01v8[cbd]
let cbs_PM3=@m.x1.XPM3.msky130_fd_pr__pfet_01v8[cbs]
let cdg_PM3=@m.x1.XPM3.msky130_fd_pr__pfet_01v8[cdg]
let cdd_PM3=@m.x1.XPM3.msky130_fd_pr__pfet_01v8[cdd]
let cds_PM3=@m.x1.XPM3.msky130_fd_pr__pfet_01v8[cds]
let csg_PM3=@m.x1.XPM3.msky130_fd_pr__pfet_01v8[csg]
let csd_PM3=@m.x1.XPM3.msky130_fd_pr__pfet_01v8[csd]
let css_PM3=@m.x1.XPM3.msky130_fd_pr__pfet_01v8[css]
let cgb_PM3=@m.x1.XPM3.msky130_fd_pr__pfet_01v8[cgb]
let cdb_PM3=@m.x1.XPM3.msky130_fd_pr__pfet_01v8[cdb]
let csb_PM3=@m.x1.XPM3.msky130_fd_pr__pfet_01v8[csb]
let cbb_PM3=@m.x1.XPM3.msky130_fd_pr__pfet_01v8[cbb]
let capbd_PM3=@m.x1.XPM3.msky130_fd_pr__pfet_01v8[capbd]
let capbs_PM3=@m.x1.XPM3.msky130_fd_pr__pfet_01v8[capbs]
let qg_PM3=@m.x1.XPM3.msky130_fd_pr__pfet_01v8[qg]
let qb_PM3=@m.x1.XPM3.msky130_fd_pr__pfet_01v8[qb]
let qs_PM3=@m.x1.XPM3.msky130_fd_pr__pfet_01v8[qs]
let qinv_PM3=@m.x1.XPM3.msky130_fd_pr__pfet_01v8[qinv]
let qdef_PM3=@m.x1.XPM3.msky130_fd_pr__pfet_01v8[qdef]
let gcrg_PM3=@m.x1.XPM3.msky130_fd_pr__pfet_01v8[gcrg]
let gtau_PM3=@m.x1.XPM3.msky130_fd_pr__pfet_01v8[gtau]

let gmbs_PM4=@m.x1.XPM4.msky130_fd_pr__pfet_01v8[gmbs]
let gm_PM4=@m.x1.XPM4.msky130_fd_pr__pfet_01v8[gm]
let gds_PM4=@m.x1.XPM4.msky130_fd_pr__pfet_01v8[gds]
let vdsat_PM4=@m.x1.XPM4.msky130_fd_pr__pfet_01v8[vdsat]
let vth_PM4=@m.x1.XPM4.msky130_fd_pr__pfet_01v8[vth]
let id_PM4=@m.x1.XPM4.msky130_fd_pr__pfet_01v8[id]
let ibd_PM4=@m.x1.XPM4.msky130_fd_pr__pfet_01v8[ibd]
let ibs_PM4=@m.x1.XPM4.msky130_fd_pr__pfet_01v8[ibs]
let gbd_PM4=@m.x1.XPM4.msky130_fd_pr__pfet_01v8[gbd]
let gbs_PM4=@m.x1.XPM4.msky130_fd_pr__pfet_01v8[gbs]
let isub_PM4=@m.x1.XPM4.msky130_fd_pr__pfet_01v8[isub]
let igidl_PM4=@m.x1.XPM4.msky130_fd_pr__pfet_01v8[igidl]
let igisl_PM4=@m.x1.XPM4.msky130_fd_pr__pfet_01v8[igisl]
let igs_PM4=@m.x1.XPM4.msky130_fd_pr__pfet_01v8[igs]
let igd_PM4=@m.x1.XPM4.msky130_fd_pr__pfet_01v8[igd]
let igb_PM4=@m.x1.XPM4.msky130_fd_pr__pfet_01v8[igb]
let igcs_PM4=@m.x1.XPM4.msky130_fd_pr__pfet_01v8[igcs]
let vbs_PM4=@m.x1.XPM4.msky130_fd_pr__pfet_01v8[vbs]
let vgs_PM4=@m.x1.XPM4.msky130_fd_pr__pfet_01v8[vgs]
let vds_PM4=@m.x1.XPM4.msky130_fd_pr__pfet_01v8[vds]
let cgg_PM4=@m.x1.XPM4.msky130_fd_pr__pfet_01v8[cgg]
let cgs_PM4=@m.x1.XPM4.msky130_fd_pr__pfet_01v8[cgs]
let cgd_PM4=@m.x1.XPM4.msky130_fd_pr__pfet_01v8[cgd]
let cbg_PM4=@m.x1.XPM4.msky130_fd_pr__pfet_01v8[cbg]
let cbd_PM4=@m.x1.XPM4.msky130_fd_pr__pfet_01v8[cbd]
let cbs_PM4=@m.x1.XPM4.msky130_fd_pr__pfet_01v8[cbs]
let cdg_PM4=@m.x1.XPM4.msky130_fd_pr__pfet_01v8[cdg]
let cdd_PM4=@m.x1.XPM4.msky130_fd_pr__pfet_01v8[cdd]
let cds_PM4=@m.x1.XPM4.msky130_fd_pr__pfet_01v8[cds]
let csg_PM4=@m.x1.XPM4.msky130_fd_pr__pfet_01v8[csg]
let csd_PM4=@m.x1.XPM4.msky130_fd_pr__pfet_01v8[csd]
let css_PM4=@m.x1.XPM4.msky130_fd_pr__pfet_01v8[css]
let cgb_PM4=@m.x1.XPM4.msky130_fd_pr__pfet_01v8[cgb]
let cdb_PM4=@m.x1.XPM4.msky130_fd_pr__pfet_01v8[cdb]
let csb_PM4=@m.x1.XPM4.msky130_fd_pr__pfet_01v8[csb]
let cbb_PM4=@m.x1.XPM4.msky130_fd_pr__pfet_01v8[cbb]
let capbd_PM4=@m.x1.XPM4.msky130_fd_pr__pfet_01v8[capbd]
let capbs_PM4=@m.x1.XPM4.msky130_fd_pr__pfet_01v8[capbs]
let qg_PM4=@m.x1.XPM4.msky130_fd_pr__pfet_01v8[qg]
let qb_PM4=@m.x1.XPM4.msky130_fd_pr__pfet_01v8[qb]
let qs_PM4=@m.x1.XPM4.msky130_fd_pr__pfet_01v8[qs]
let qinv_PM4=@m.x1.XPM4.msky130_fd_pr__pfet_01v8[qinv]
let qdef_PM4=@m.x1.XPM4.msky130_fd_pr__pfet_01v8[qdef]
let gcrg_PM4=@m.x1.XPM4.msky130_fd_pr__pfet_01v8[gcrg]
let gtau_PM4=@m.x1.XPM4.msky130_fd_pr__pfet_01v8[gtau]

let gmbs_PM5=@m.x1.XPM5.msky130_fd_pr__pfet_01v8[gmbs]
let gm_PM5=@m.x1.XPM5.msky130_fd_pr__pfet_01v8[gm]
let gds_PM5=@m.x1.XPM5.msky130_fd_pr__pfet_01v8[gds]
let vdsat_PM5=@m.x1.XPM5.msky130_fd_pr__pfet_01v8[vdsat]
let vth_PM5=@m.x1.XPM5.msky130_fd_pr__pfet_01v8[vth]
let id_PM5=@m.x1.XPM5.msky130_fd_pr__pfet_01v8[id]
let ibd_PM5=@m.x1.XPM5.msky130_fd_pr__pfet_01v8[ibd]
let ibs_PM5=@m.x1.XPM5.msky130_fd_pr__pfet_01v8[ibs]
let gbd_PM5=@m.x1.XPM5.msky130_fd_pr__pfet_01v8[gbd]
let gbs_PM5=@m.x1.XPM5.msky130_fd_pr__pfet_01v8[gbs]
let isub_PM5=@m.x1.XPM5.msky130_fd_pr__pfet_01v8[isub]
let igidl_PM5=@m.x1.XPM5.msky130_fd_pr__pfet_01v8[igidl]
let igisl_PM5=@m.x1.XPM5.msky130_fd_pr__pfet_01v8[igisl]
let igs_PM5=@m.x1.XPM5.msky130_fd_pr__pfet_01v8[igs]
let igd_PM5=@m.x1.XPM5.msky130_fd_pr__pfet_01v8[igd]
let igb_PM5=@m.x1.XPM5.msky130_fd_pr__pfet_01v8[igb]
let igcs_PM5=@m.x1.XPM5.msky130_fd_pr__pfet_01v8[igcs]
let vbs_PM5=@m.x1.XPM5.msky130_fd_pr__pfet_01v8[vbs]
let vgs_PM5=@m.x1.XPM5.msky130_fd_pr__pfet_01v8[vgs]
let vds_PM5=@m.x1.XPM5.msky130_fd_pr__pfet_01v8[vds]
let cgg_PM5=@m.x1.XPM5.msky130_fd_pr__pfet_01v8[cgg]
let cgs_PM5=@m.x1.XPM5.msky130_fd_pr__pfet_01v8[cgs]
let cgd_PM5=@m.x1.XPM5.msky130_fd_pr__pfet_01v8[cgd]
let cbg_PM5=@m.x1.XPM5.msky130_fd_pr__pfet_01v8[cbg]
let cbd_PM5=@m.x1.XPM5.msky130_fd_pr__pfet_01v8[cbd]
let cbs_PM5=@m.x1.XPM5.msky130_fd_pr__pfet_01v8[cbs]
let cdg_PM5=@m.x1.XPM5.msky130_fd_pr__pfet_01v8[cdg]
let cdd_PM5=@m.x1.XPM5.msky130_fd_pr__pfet_01v8[cdd]
let cds_PM5=@m.x1.XPM5.msky130_fd_pr__pfet_01v8[cds]
let csg_PM5=@m.x1.XPM5.msky130_fd_pr__pfet_01v8[csg]
let csd_PM5=@m.x1.XPM5.msky130_fd_pr__pfet_01v8[csd]
let css_PM5=@m.x1.XPM5.msky130_fd_pr__pfet_01v8[css]
let cgb_PM5=@m.x1.XPM5.msky130_fd_pr__pfet_01v8[cgb]
let cdb_PM5=@m.x1.XPM5.msky130_fd_pr__pfet_01v8[cdb]
let csb_PM5=@m.x1.XPM5.msky130_fd_pr__pfet_01v8[csb]
let cbb_PM5=@m.x1.XPM5.msky130_fd_pr__pfet_01v8[cbb]
let capbd_PM5=@m.x1.XPM5.msky130_fd_pr__pfet_01v8[capbd]
let capbs_PM5=@m.x1.XPM5.msky130_fd_pr__pfet_01v8[capbs]
let qg_PM5=@m.x1.XPM5.msky130_fd_pr__pfet_01v8[qg]
let qb_PM5=@m.x1.XPM5.msky130_fd_pr__pfet_01v8[qb]
let qs_PM5=@m.x1.XPM5.msky130_fd_pr__pfet_01v8[qs]
let qinv_PM5=@m.x1.XPM5.msky130_fd_pr__pfet_01v8[qinv]
let qdef_PM5=@m.x1.XPM5.msky130_fd_pr__pfet_01v8[qdef]
let gcrg_PM5=@m.x1.XPM5.msky130_fd_pr__pfet_01v8[gcrg]
let gtau_PM5=@m.x1.XPM5.msky130_fd_pr__pfet_01v8[gtau]

let gmbs_PM6=@m.x1.XPM6.msky130_fd_pr__pfet_01v8[gmbs]
let gm_PM6=@m.x1.XPM6.msky130_fd_pr__pfet_01v8[gm]
let gds_PM6=@m.x1.XPM6.msky130_fd_pr__pfet_01v8[gds]
let vdsat_PM6=@m.x1.XPM6.msky130_fd_pr__pfet_01v8[vdsat]
let vth_PM6=@m.x1.XPM6.msky130_fd_pr__pfet_01v8[vth]
let id_PM6=@m.x1.XPM6.msky130_fd_pr__pfet_01v8[id]
let ibd_PM6=@m.x1.XPM6.msky130_fd_pr__pfet_01v8[ibd]
let ibs_PM6=@m.x1.XPM6.msky130_fd_pr__pfet_01v8[ibs]
let gbd_PM6=@m.x1.XPM6.msky130_fd_pr__pfet_01v8[gbd]
let gbs_PM6=@m.x1.XPM6.msky130_fd_pr__pfet_01v8[gbs]
let isub_PM6=@m.x1.XPM6.msky130_fd_pr__pfet_01v8[isub]
let igidl_PM6=@m.x1.XPM6.msky130_fd_pr__pfet_01v8[igidl]
let igisl_PM6=@m.x1.XPM6.msky130_fd_pr__pfet_01v8[igisl]
let igs_PM6=@m.x1.XPM6.msky130_fd_pr__pfet_01v8[igs]
let igd_PM6=@m.x1.XPM6.msky130_fd_pr__pfet_01v8[igd]
let igb_PM6=@m.x1.XPM6.msky130_fd_pr__pfet_01v8[igb]
let igcs_PM6=@m.x1.XPM6.msky130_fd_pr__pfet_01v8[igcs]
let vbs_PM6=@m.x1.XPM6.msky130_fd_pr__pfet_01v8[vbs]
let vgs_PM6=@m.x1.XPM6.msky130_fd_pr__pfet_01v8[vgs]
let vds_PM6=@m.x1.XPM6.msky130_fd_pr__pfet_01v8[vds]
let cgg_PM6=@m.x1.XPM6.msky130_fd_pr__pfet_01v8[cgg]
let cgs_PM6=@m.x1.XPM6.msky130_fd_pr__pfet_01v8[cgs]
let cgd_PM6=@m.x1.XPM6.msky130_fd_pr__pfet_01v8[cgd]
let cbg_PM6=@m.x1.XPM6.msky130_fd_pr__pfet_01v8[cbg]
let cbd_PM6=@m.x1.XPM6.msky130_fd_pr__pfet_01v8[cbd]
let cbs_PM6=@m.x1.XPM6.msky130_fd_pr__pfet_01v8[cbs]
let cdg_PM6=@m.x1.XPM6.msky130_fd_pr__pfet_01v8[cdg]
let cdd_PM6=@m.x1.XPM6.msky130_fd_pr__pfet_01v8[cdd]
let cds_PM6=@m.x1.XPM6.msky130_fd_pr__pfet_01v8[cds]
let csg_PM6=@m.x1.XPM6.msky130_fd_pr__pfet_01v8[csg]
let csd_PM6=@m.x1.XPM6.msky130_fd_pr__pfet_01v8[csd]
let css_PM6=@m.x1.XPM6.msky130_fd_pr__pfet_01v8[css]
let cgb_PM6=@m.x1.XPM6.msky130_fd_pr__pfet_01v8[cgb]
let cdb_PM6=@m.x1.XPM6.msky130_fd_pr__pfet_01v8[cdb]
let csb_PM6=@m.x1.XPM6.msky130_fd_pr__pfet_01v8[csb]
let cbb_PM6=@m.x1.XPM6.msky130_fd_pr__pfet_01v8[cbb]
let capbd_PM6=@m.x1.XPM6.msky130_fd_pr__pfet_01v8[capbd]
let capbs_PM6=@m.x1.XPM6.msky130_fd_pr__pfet_01v8[capbs]
let qg_PM6=@m.x1.XPM6.msky130_fd_pr__pfet_01v8[qg]
let qb_PM6=@m.x1.XPM6.msky130_fd_pr__pfet_01v8[qb]
let qs_PM6=@m.x1.XPM6.msky130_fd_pr__pfet_01v8[qs]
let qinv_PM6=@m.x1.XPM6.msky130_fd_pr__pfet_01v8[qinv]
let qdef_PM6=@m.x1.XPM6.msky130_fd_pr__pfet_01v8[qdef]
let gcrg_PM6=@m.x1.XPM6.msky130_fd_pr__pfet_01v8[gcrg]
let gtau_PM6=@m.x1.XPM6.msky130_fd_pr__pfet_01v8[gtau]

let gmbs_PM7=@m.x1.XPM7.msky130_fd_pr__pfet_01v8[gmbs]
let gm_PM7=@m.x1.XPM7.msky130_fd_pr__pfet_01v8[gm]
let gds_PM7=@m.x1.XPM7.msky130_fd_pr__pfet_01v8[gds]
let vdsat_PM7=@m.x1.XPM7.msky130_fd_pr__pfet_01v8[vdsat]
let vth_PM7=@m.x1.XPM7.msky130_fd_pr__pfet_01v8[vth]
let id_PM7=@m.x1.XPM7.msky130_fd_pr__pfet_01v8[id]
let ibd_PM7=@m.x1.XPM7.msky130_fd_pr__pfet_01v8[ibd]
let ibs_PM7=@m.x1.XPM7.msky130_fd_pr__pfet_01v8[ibs]
let gbd_PM7=@m.x1.XPM7.msky130_fd_pr__pfet_01v8[gbd]
let gbs_PM7=@m.x1.XPM7.msky130_fd_pr__pfet_01v8[gbs]
let isub_PM7=@m.x1.XPM7.msky130_fd_pr__pfet_01v8[isub]
let igidl_PM7=@m.x1.XPM7.msky130_fd_pr__pfet_01v8[igidl]
let igisl_PM7=@m.x1.XPM7.msky130_fd_pr__pfet_01v8[igisl]
let igs_PM7=@m.x1.XPM7.msky130_fd_pr__pfet_01v8[igs]
let igd_PM7=@m.x1.XPM7.msky130_fd_pr__pfet_01v8[igd]
let igb_PM7=@m.x1.XPM7.msky130_fd_pr__pfet_01v8[igb]
let igcs_PM7=@m.x1.XPM7.msky130_fd_pr__pfet_01v8[igcs]
let vbs_PM7=@m.x1.XPM7.msky130_fd_pr__pfet_01v8[vbs]
let vgs_PM7=@m.x1.XPM7.msky130_fd_pr__pfet_01v8[vgs]
let vds_PM7=@m.x1.XPM7.msky130_fd_pr__pfet_01v8[vds]
let cgg_PM7=@m.x1.XPM7.msky130_fd_pr__pfet_01v8[cgg]
let cgs_PM7=@m.x1.XPM7.msky130_fd_pr__pfet_01v8[cgs]
let cgd_PM7=@m.x1.XPM7.msky130_fd_pr__pfet_01v8[cgd]
let cbg_PM7=@m.x1.XPM7.msky130_fd_pr__pfet_01v8[cbg]
let cbd_PM7=@m.x1.XPM7.msky130_fd_pr__pfet_01v8[cbd]
let cbs_PM7=@m.x1.XPM7.msky130_fd_pr__pfet_01v8[cbs]
let cdg_PM7=@m.x1.XPM7.msky130_fd_pr__pfet_01v8[cdg]
let cdd_PM7=@m.x1.XPM7.msky130_fd_pr__pfet_01v8[cdd]
let cds_PM7=@m.x1.XPM7.msky130_fd_pr__pfet_01v8[cds]
let csg_PM7=@m.x1.XPM7.msky130_fd_pr__pfet_01v8[csg]
let csd_PM7=@m.x1.XPM7.msky130_fd_pr__pfet_01v8[csd]
let css_PM7=@m.x1.XPM7.msky130_fd_pr__pfet_01v8[css]
let cgb_PM7=@m.x1.XPM7.msky130_fd_pr__pfet_01v8[cgb]
let cdb_PM7=@m.x1.XPM7.msky130_fd_pr__pfet_01v8[cdb]
let csb_PM7=@m.x1.XPM7.msky130_fd_pr__pfet_01v8[csb]
let cbb_PM7=@m.x1.XPM7.msky130_fd_pr__pfet_01v8[cbb]
let capbd_PM7=@m.x1.XPM7.msky130_fd_pr__pfet_01v8[capbd]
let capbs_PM7=@m.x1.XPM7.msky130_fd_pr__pfet_01v8[capbs]
let qg_PM7=@m.x1.XPM7.msky130_fd_pr__pfet_01v8[qg]
let qb_PM7=@m.x1.XPM7.msky130_fd_pr__pfet_01v8[qb]
let qs_PM7=@m.x1.XPM7.msky130_fd_pr__pfet_01v8[qs]
let qinv_PM7=@m.x1.XPM7.msky130_fd_pr__pfet_01v8[qinv]
let qdef_PM7=@m.x1.XPM7.msky130_fd_pr__pfet_01v8[qdef]
let gcrg_PM7=@m.x1.XPM7.msky130_fd_pr__pfet_01v8[gcrg]
let gtau_PM7=@m.x1.XPM7.msky130_fd_pr__pfet_01v8[gtau]

let gmbs_PM8=@m.x1.XPM8.msky130_fd_pr__pfet_01v8[gmbs]
let gm_PM8=@m.x1.XPM8.msky130_fd_pr__pfet_01v8[gm]
let gds_PM8=@m.x1.XPM8.msky130_fd_pr__pfet_01v8[gds]
let vdsat_PM8=@m.x1.XPM8.msky130_fd_pr__pfet_01v8[vdsat]
let vth_PM8=@m.x1.XPM8.msky130_fd_pr__pfet_01v8[vth]
let id_PM8=@m.x1.XPM8.msky130_fd_pr__pfet_01v8[id]
let ibd_PM8=@m.x1.XPM8.msky130_fd_pr__pfet_01v8[ibd]
let ibs_PM8=@m.x1.XPM8.msky130_fd_pr__pfet_01v8[ibs]
let gbd_PM8=@m.x1.XPM8.msky130_fd_pr__pfet_01v8[gbd]
let gbs_PM8=@m.x1.XPM8.msky130_fd_pr__pfet_01v8[gbs]
let isub_PM8=@m.x1.XPM8.msky130_fd_pr__pfet_01v8[isub]
let igidl_PM8=@m.x1.XPM8.msky130_fd_pr__pfet_01v8[igidl]
let igisl_PM8=@m.x1.XPM8.msky130_fd_pr__pfet_01v8[igisl]
let igs_PM8=@m.x1.XPM8.msky130_fd_pr__pfet_01v8[igs]
let igd_PM8=@m.x1.XPM8.msky130_fd_pr__pfet_01v8[igd]
let igb_PM8=@m.x1.XPM8.msky130_fd_pr__pfet_01v8[igb]
let igcs_PM8=@m.x1.XPM8.msky130_fd_pr__pfet_01v8[igcs]
let vbs_PM8=@m.x1.XPM8.msky130_fd_pr__pfet_01v8[vbs]
let vgs_PM8=@m.x1.XPM8.msky130_fd_pr__pfet_01v8[vgs]
let vds_PM8=@m.x1.XPM8.msky130_fd_pr__pfet_01v8[vds]
let cgg_PM8=@m.x1.XPM8.msky130_fd_pr__pfet_01v8[cgg]
let cgs_PM8=@m.x1.XPM8.msky130_fd_pr__pfet_01v8[cgs]
let cgd_PM8=@m.x1.XPM8.msky130_fd_pr__pfet_01v8[cgd]
let cbg_PM8=@m.x1.XPM8.msky130_fd_pr__pfet_01v8[cbg]
let cbd_PM8=@m.x1.XPM8.msky130_fd_pr__pfet_01v8[cbd]
let cbs_PM8=@m.x1.XPM8.msky130_fd_pr__pfet_01v8[cbs]
let cdg_PM8=@m.x1.XPM8.msky130_fd_pr__pfet_01v8[cdg]
let cdd_PM8=@m.x1.XPM8.msky130_fd_pr__pfet_01v8[cdd]
let cds_PM8=@m.x1.XPM8.msky130_fd_pr__pfet_01v8[cds]
let csg_PM8=@m.x1.XPM8.msky130_fd_pr__pfet_01v8[csg]
let csd_PM8=@m.x1.XPM8.msky130_fd_pr__pfet_01v8[csd]
let css_PM8=@m.x1.XPM8.msky130_fd_pr__pfet_01v8[css]
let cgb_PM8=@m.x1.XPM8.msky130_fd_pr__pfet_01v8[cgb]
let cdb_PM8=@m.x1.XPM8.msky130_fd_pr__pfet_01v8[cdb]
let csb_PM8=@m.x1.XPM8.msky130_fd_pr__pfet_01v8[csb]
let cbb_PM8=@m.x1.XPM8.msky130_fd_pr__pfet_01v8[cbb]
let capbd_PM8=@m.x1.XPM8.msky130_fd_pr__pfet_01v8[capbd]
let capbs_PM8=@m.x1.XPM8.msky130_fd_pr__pfet_01v8[capbs]
let qg_PM8=@m.x1.XPM8.msky130_fd_pr__pfet_01v8[qg]
let qb_PM8=@m.x1.XPM8.msky130_fd_pr__pfet_01v8[qb]
let qs_PM8=@m.x1.XPM8.msky130_fd_pr__pfet_01v8[qs]
let qinv_PM8=@m.x1.XPM8.msky130_fd_pr__pfet_01v8[qinv]
let qdef_PM8=@m.x1.XPM8.msky130_fd_pr__pfet_01v8[qdef]
let gcrg_PM8=@m.x1.XPM8.msky130_fd_pr__pfet_01v8[gcrg]
let gtau_PM8=@m.x1.XPM8.msky130_fd_pr__pfet_01v8[gtau]

let gmbs_PM9=@m.x1.XPM9.msky130_fd_pr__pfet_01v8[gmbs]
let gm_PM9=@m.x1.XPM9.msky130_fd_pr__pfet_01v8[gm]
let gds_PM9=@m.x1.XPM9.msky130_fd_pr__pfet_01v8[gds]
let vdsat_PM9=@m.x1.XPM9.msky130_fd_pr__pfet_01v8[vdsat]
let vth_PM9=@m.x1.XPM9.msky130_fd_pr__pfet_01v8[vth]
let id_PM9=@m.x1.XPM9.msky130_fd_pr__pfet_01v8[id]
let ibd_PM9=@m.x1.XPM9.msky130_fd_pr__pfet_01v8[ibd]
let ibs_PM9=@m.x1.XPM9.msky130_fd_pr__pfet_01v8[ibs]
let gbd_PM9=@m.x1.XPM9.msky130_fd_pr__pfet_01v8[gbd]
let gbs_PM9=@m.x1.XPM9.msky130_fd_pr__pfet_01v8[gbs]
let isub_PM9=@m.x1.XPM9.msky130_fd_pr__pfet_01v8[isub]
let igidl_PM9=@m.x1.XPM9.msky130_fd_pr__pfet_01v8[igidl]
let igisl_PM9=@m.x1.XPM9.msky130_fd_pr__pfet_01v8[igisl]
let igs_PM9=@m.x1.XPM9.msky130_fd_pr__pfet_01v8[igs]
let igd_PM9=@m.x1.XPM9.msky130_fd_pr__pfet_01v8[igd]
let igb_PM9=@m.x1.XPM9.msky130_fd_pr__pfet_01v8[igb]
let igcs_PM9=@m.x1.XPM9.msky130_fd_pr__pfet_01v8[igcs]
let vbs_PM9=@m.x1.XPM9.msky130_fd_pr__pfet_01v8[vbs]
let vgs_PM9=@m.x1.XPM9.msky130_fd_pr__pfet_01v8[vgs]
let vds_PM9=@m.x1.XPM9.msky130_fd_pr__pfet_01v8[vds]
let cgg_PM9=@m.x1.XPM9.msky130_fd_pr__pfet_01v8[cgg]
let cgs_PM9=@m.x1.XPM9.msky130_fd_pr__pfet_01v8[cgs]
let cgd_PM9=@m.x1.XPM9.msky130_fd_pr__pfet_01v8[cgd]
let cbg_PM9=@m.x1.XPM9.msky130_fd_pr__pfet_01v8[cbg]
let cbd_PM9=@m.x1.XPM9.msky130_fd_pr__pfet_01v8[cbd]
let cbs_PM9=@m.x1.XPM9.msky130_fd_pr__pfet_01v8[cbs]
let cdg_PM9=@m.x1.XPM9.msky130_fd_pr__pfet_01v8[cdg]
let cdd_PM9=@m.x1.XPM9.msky130_fd_pr__pfet_01v8[cdd]
let cds_PM9=@m.x1.XPM9.msky130_fd_pr__pfet_01v8[cds]
let csg_PM9=@m.x1.XPM9.msky130_fd_pr__pfet_01v8[csg]
let csd_PM9=@m.x1.XPM9.msky130_fd_pr__pfet_01v8[csd]
let css_PM9=@m.x1.XPM9.msky130_fd_pr__pfet_01v8[css]
let cgb_PM9=@m.x1.XPM9.msky130_fd_pr__pfet_01v8[cgb]
let cdb_PM9=@m.x1.XPM9.msky130_fd_pr__pfet_01v8[cdb]
let csb_PM9=@m.x1.XPM9.msky130_fd_pr__pfet_01v8[csb]
let cbb_PM9=@m.x1.XPM9.msky130_fd_pr__pfet_01v8[cbb]
let capbd_PM9=@m.x1.XPM9.msky130_fd_pr__pfet_01v8[capbd]
let capbs_PM9=@m.x1.XPM9.msky130_fd_pr__pfet_01v8[capbs]
let qg_PM9=@m.x1.XPM9.msky130_fd_pr__pfet_01v8[qg]
let qb_PM9=@m.x1.XPM9.msky130_fd_pr__pfet_01v8[qb]
let qs_PM9=@m.x1.XPM9.msky130_fd_pr__pfet_01v8[qs]
let qinv_PM9=@m.x1.XPM9.msky130_fd_pr__pfet_01v8[qinv]
let qdef_PM9=@m.x1.XPM9.msky130_fd_pr__pfet_01v8[qdef]
let gcrg_PM9=@m.x1.XPM9.msky130_fd_pr__pfet_01v8[gcrg]
let gtau_PM9=@m.x1.XPM9.msky130_fd_pr__pfet_01v8[gtau]

let dc_Ib=@Ib[dc]
let acmag_Ib=@Ib[acmag]
let acphase_Ib=@Ib[acphase]
let acreal_Ib=@Ib[acreal]
let acimag_Ib=@Ib[acimag]
let v_Ib=@Ib[v]
let p_Ib=@Ib[p]
let current_Ib=@Ib[current]

let capacitance_C0=@c.x1.XC0.c1[capacitance]
let cap_C0=@c.x1.XC0.c1[cap]
let c_C0=@c.x1.XC0.c1[c]
let ic_C0=@c.x1.XC0.c1[ic]
let temp_C0=@c.x1.XC0.c1[temp]
let dtemp_C0=@c.x1.XC0.c1[dtemp]
let w_C0=@c.x1.XC0.c1[w]
let l_C0=@c.x1.XC0.c1[l]
let m_C0=@c.x1.XC0.c1[m]
let scale_C0=@c.x1.XC0.c1[scale]
let i_C0=@c.x1.XC0.c1[i]
let p_C0=@c.x1.XC0.c1[p]
let sens_dc_C0=@c.x1.XC0.c1[sens_dc]
let sens_real_C0=@c.x1.XC0.c1[sens_real]
let sens_imag_C0=@c.x1.XC0.c1[sens_imag]
let sens_mag_C0=@c.x1.XC0.c1[sens_mag]
let sens_ph_C0=@c.x1.XC0.c1[sens_ph]
let sens_cplx_C0=@c.x1.XC0.c1[sens_cplx]

let capacitance_C1=@c.x1.XC1.c1[capacitance]
let cap_C1=@c.x1.XC1.c1[cap]
let c_C1=@c.x1.XC1.c1[c]
let ic_C1=@c.x1.XC1.c1[ic]
let temp_C1=@c.x1.XC1.c1[temp]
let dtemp_C1=@c.x1.XC1.c1[dtemp]
let w_C1=@c.x1.XC1.c1[w]
let l_C1=@c.x1.XC1.c1[l]
let m_C1=@c.x1.XC1.c1[m]
let scale_C1=@c.x1.XC1.c1[scale]
let i_C1=@c.x1.XC1.c1[i]
let p_C1=@c.x1.XC1.c1[p]
let sens_dc_C1=@c.x1.XC1.c1[sens_dc]
let sens_real_C1=@c.x1.XC1.c1[sens_real]
let sens_imag_C1=@c.x1.XC1.c1[sens_imag]
let sens_mag_C1=@c.x1.XC1.c1[sens_mag]
let sens_ph_C1=@c.x1.XC1.c1[sens_ph]
let sens_cplx_C1=@c.x1.XC1.c1[sens_cplx]

let capacitance_C4=@c.x1.XC4.c1[capacitance]
let cap_C4=@c.x1.XC4.c1[cap]
let c_C4=@c.x1.XC4.c1[c]
let ic_C4=@c.x1.XC4.c1[ic]
let temp_C4=@c.x1.XC4.c1[temp]
let dtemp_C4=@c.x1.XC4.c1[dtemp]
let w_C4=@c.x1.XC4.c1[w]
let l_C4=@c.x1.XC4.c1[l]
let m_C4=@c.x1.XC4.c1[m]
let scale_C4=@c.x1.XC4.c1[scale]
let i_C4=@c.x1.XC4.c1[i]
let p_C4=@c.x1.XC4.c1[p]
let sens_dc_C4=@c.x1.XC4.c1[sens_dc]
let sens_real_C4=@c.x1.XC4.c1[sens_real]
let sens_imag_C4=@c.x1.XC4.c1[sens_imag]
let sens_mag_C4=@c.x1.XC4.c1[sens_mag]
let sens_ph_C4=@c.x1.XC4.c1[sens_ph]
let sens_cplx_C4=@c.x1.XC4.c1[sens_cplx]

let capacitance_CL=@c.XCL.c1[capacitance]
let cap_CL=@c.XCL.c1[cap]
let c_CL=@c.XCL.c1[c]
let ic_CL=@c.XCL.c1[ic]
let temp_CL=@c.XCL.c1[temp]
let dtemp_CL=@c.XCL.c1[dtemp]
let w_CL=@c.XCL.c1[w]
let l_CL=@c.XCL.c1[l]
let m_CL=@c.XCL.c1[m]
let scale_CL=@c.XCL.c1[scale]
let i_CL=@c.XCL.c1[i]
let p_CL=@c.XCL.c1[p]
let sens_dc_CL=@c.XCL.c1[sens_dc]
let sens_real_CL=@c.XCL.c1[sens_real]
let sens_imag_CL=@c.XCL.c1[sens_imag]
let sens_mag_CL=@c.XCL.c1[sens_mag]
let sens_ph_CL=@c.XCL.c1[sens_ph]
let sens_cplx_CL=@c.XCL.c1[sens_cplx]

write ldo_2_op gmbs_NM0 gm_NM0 gds_NM0 vdsat_NM0 vth_NM0 id_NM0 ibd_NM0 ibs_NM0 gbd_NM0 gbs_NM0 isub_NM0 igidl_NM0 igisl_NM0 igs_NM0 igd_NM0 igb_NM0 igcs_NM0 vbs_NM0 vgs_NM0 vds_NM0 cgg_NM0 cgs_NM0 cgd_NM0 cbg_NM0 cbd_NM0 cbs_NM0 cdg_NM0 cdd_NM0 cds_NM0 csg_NM0 csd_NM0 css_NM0 cgb_NM0 cdb_NM0 csb_NM0 cbb_NM0 capbd_NM0 capbs_NM0 qg_NM0 qb_NM0 qs_NM0 qinv_NM0 qdef_NM0 gcrg_NM0 gtau_NM0 gmbs_NM1 gm_NM1 gds_NM1 vdsat_NM1 vth_NM1 id_NM1 ibd_NM1 ibs_NM1 gbd_NM1 gbs_NM1 isub_NM1 igidl_NM1 igisl_NM1 igs_NM1 igd_NM1 igb_NM1 igcs_NM1 vbs_NM1 vgs_NM1 vds_NM1 cgg_NM1 cgs_NM1 cgd_NM1 cbg_NM1 cbd_NM1 cbs_NM1 cdg_NM1 cdd_NM1 cds_NM1 csg_NM1 csd_NM1 css_NM1 cgb_NM1 cdb_NM1 csb_NM1 cbb_NM1 capbd_NM1 capbs_NM1 qg_NM1 qb_NM1 qs_NM1 qinv_NM1 qdef_NM1 gcrg_NM1 gtau_NM1 gmbs_NM2 gm_NM2 gds_NM2 vdsat_NM2 vth_NM2 id_NM2 ibd_NM2 ibs_NM2 gbd_NM2 gbs_NM2 isub_NM2 igidl_NM2 igisl_NM2 igs_NM2 igd_NM2 igb_NM2 igcs_NM2 vbs_NM2 vgs_NM2 vds_NM2 cgg_NM2 cgs_NM2 cgd_NM2 cbg_NM2 cbd_NM2 cbs_NM2 cdg_NM2 cdd_NM2 cds_NM2 csg_NM2 csd_NM2 css_NM2 cgb_NM2 cdb_NM2 csb_NM2 cbb_NM2 capbd_NM2 capbs_NM2 qg_NM2 qb_NM2 qs_NM2 qinv_NM2 qdef_NM2 gcrg_NM2 gtau_NM2 gmbs_NM3 gm_NM3 gds_NM3 vdsat_NM3 vth_NM3 id_NM3 ibd_NM3 ibs_NM3 gbd_NM3 gbs_NM3 isub_NM3 igidl_NM3 igisl_NM3 igs_NM3 igd_NM3 igb_NM3 igcs_NM3 vbs_NM3 vgs_NM3 vds_NM3 cgg_NM3 cgs_NM3 cgd_NM3 cbg_NM3 cbd_NM3 cbs_NM3 cdg_NM3 cdd_NM3 cds_NM3 csg_NM3 csd_NM3 css_NM3 cgb_NM3 cdb_NM3 csb_NM3 cbb_NM3 capbd_NM3 capbs_NM3 qg_NM3 qb_NM3 qs_NM3 qinv_NM3 qdef_NM3 gcrg_NM3 gtau_NM3 gmbs_NM4 gm_NM4 gds_NM4 vdsat_NM4 vth_NM4 id_NM4 ibd_NM4 ibs_NM4 gbd_NM4 gbs_NM4 isub_NM4 igidl_NM4 igisl_NM4 igs_NM4 igd_NM4 igb_NM4 igcs_NM4 vbs_NM4 vgs_NM4 vds_NM4 cgg_NM4 cgs_NM4 cgd_NM4 cbg_NM4 cbd_NM4 cbs_NM4 cdg_NM4 cdd_NM4 cds_NM4 csg_NM4 csd_NM4 css_NM4 cgb_NM4 cdb_NM4 csb_NM4 cbb_NM4 capbd_NM4 capbs_NM4 qg_NM4 qb_NM4 qs_NM4 qinv_NM4 qdef_NM4 gcrg_NM4 gtau_NM4 gmbs_NM6 gm_NM6 gds_NM6 vdsat_NM6 vth_NM6 id_NM6 ibd_NM6 ibs_NM6 gbd_NM6 gbs_NM6 isub_NM6 igidl_NM6 igisl_NM6 igs_NM6 igd_NM6 igb_NM6 igcs_NM6 vbs_NM6 vgs_NM6 vds_NM6 cgg_NM6 cgs_NM6 cgd_NM6 cbg_NM6 cbd_NM6 cbs_NM6 cdg_NM6 cdd_NM6 cds_NM6 csg_NM6 csd_NM6 css_NM6 cgb_NM6 cdb_NM6 csb_NM6 cbb_NM6 capbd_NM6 capbs_NM6 qg_NM6 qb_NM6 qs_NM6 qinv_NM6 qdef_NM6 gcrg_NM6 gtau_NM6 gmbs_NM7 gm_NM7 gds_NM7 vdsat_NM7 vth_NM7 id_NM7 ibd_NM7 ibs_NM7 gbd_NM7 gbs_NM7 isub_NM7 igidl_NM7 igisl_NM7 igs_NM7 igd_NM7 igb_NM7 igcs_NM7 vbs_NM7 vgs_NM7 vds_NM7 cgg_NM7 cgs_NM7 cgd_NM7 cbg_NM7 cbd_NM7 cbs_NM7 cdg_NM7 cdd_NM7 cds_NM7 csg_NM7 csd_NM7 css_NM7 cgb_NM7 cdb_NM7 csb_NM7 cbb_NM7 capbd_NM7 capbs_NM7 qg_NM7 qb_NM7 qs_NM7 qinv_NM7 qdef_NM7 gcrg_NM7 gtau_NM7 gmbs_NM8 gm_NM8 gds_NM8 vdsat_NM8 vth_NM8 id_NM8 ibd_NM8 ibs_NM8 gbd_NM8 gbs_NM8 isub_NM8 igidl_NM8 igisl_NM8 igs_NM8 igd_NM8 igb_NM8 igcs_NM8 vbs_NM8 vgs_NM8 vds_NM8 cgg_NM8 cgs_NM8 cgd_NM8 cbg_NM8 cbd_NM8 cbs_NM8 cdg_NM8 cdd_NM8 cds_NM8 csg_NM8 csd_NM8 css_NM8 cgb_NM8 cdb_NM8 csb_NM8 cbb_NM8 capbd_NM8 capbs_NM8 qg_NM8 qb_NM8 qs_NM8 qinv_NM8 qdef_NM8 gcrg_NM8 gtau_NM8 gmbs_NM9 gm_NM9 gds_NM9 vdsat_NM9 vth_NM9 id_NM9 ibd_NM9 ibs_NM9 gbd_NM9 gbs_NM9 isub_NM9 igidl_NM9 igisl_NM9 igs_NM9 igd_NM9 igb_NM9 igcs_NM9 vbs_NM9 vgs_NM9 vds_NM9 cgg_NM9 cgs_NM9 cgd_NM9 cbg_NM9 cbd_NM9 cbs_NM9 cdg_NM9 cdd_NM9 cds_NM9 csg_NM9 csd_NM9 css_NM9 cgb_NM9 cdb_NM9 csb_NM9 cbb_NM9 capbd_NM9 capbs_NM9 qg_NM9 qb_NM9 qs_NM9 qinv_NM9 qdef_NM9 gcrg_NM9 gtau_NM9 gmbs_NM10 gm_NM10 gds_NM10 vdsat_NM10 vth_NM10 id_NM10 ibd_NM10 ibs_NM10 gbd_NM10 gbs_NM10 isub_NM10 igidl_NM10 igisl_NM10 igs_NM10 igd_NM10 igb_NM10 igcs_NM10 vbs_NM10 vgs_NM10 vds_NM10 cgg_NM10 cgs_NM10 cgd_NM10 cbg_NM10 cbd_NM10 cbs_NM10 cdg_NM10 cdd_NM10 cds_NM10 csg_NM10 csd_NM10 css_NM10 cgb_NM10 cdb_NM10 csb_NM10 cbb_NM10 capbd_NM10 capbs_NM10 qg_NM10 qb_NM10 qs_NM10 qinv_NM10 qdef_NM10 gcrg_NM10 gtau_NM10 gmbs_PM0 gm_PM0 gds_PM0 vdsat_PM0 vth_PM0 id_PM0 ibd_PM0 ibs_PM0 gbd_PM0 gbs_PM0 isub_PM0 igidl_PM0 igisl_PM0 igs_PM0 igd_PM0 igb_PM0 igcs_PM0 vbs_PM0 vgs_PM0 vds_PM0 cgg_PM0 cgs_PM0 cgd_PM0 cbg_PM0 cbd_PM0 cbs_PM0 cdg_PM0 cdd_PM0 cds_PM0 csg_PM0 csd_PM0 css_PM0 cgb_PM0 cdb_PM0 csb_PM0 cbb_PM0 capbd_PM0 capbs_PM0 qg_PM0 qb_PM0 qs_PM0 qinv_PM0 qdef_PM0 gcrg_PM0 gtau_PM0 gmbs_PM1 gm_PM1 gds_PM1 vdsat_PM1 vth_PM1 id_PM1 ibd_PM1 ibs_PM1 gbd_PM1 gbs_PM1 isub_PM1 igidl_PM1 igisl_PM1 igs_PM1 igd_PM1 igb_PM1 igcs_PM1 vbs_PM1 vgs_PM1 vds_PM1 cgg_PM1 cgs_PM1 cgd_PM1 cbg_PM1 cbd_PM1 cbs_PM1 cdg_PM1 cdd_PM1 cds_PM1 csg_PM1 csd_PM1 css_PM1 cgb_PM1 cdb_PM1 csb_PM1 cbb_PM1 capbd_PM1 capbs_PM1 qg_PM1 qb_PM1 qs_PM1 qinv_PM1 qdef_PM1 gcrg_PM1 gtau_PM1 gmbs_PM2 gm_PM2 gds_PM2 vdsat_PM2 vth_PM2 id_PM2 ibd_PM2 ibs_PM2 gbd_PM2 gbs_PM2 isub_PM2 igidl_PM2 igisl_PM2 igs_PM2 igd_PM2 igb_PM2 igcs_PM2 vbs_PM2 vgs_PM2 vds_PM2 cgg_PM2 cgs_PM2 cgd_PM2 cbg_PM2 cbd_PM2 cbs_PM2 cdg_PM2 cdd_PM2 cds_PM2 csg_PM2 csd_PM2 css_PM2 cgb_PM2 cdb_PM2 csb_PM2 cbb_PM2 capbd_PM2 capbs_PM2 qg_PM2 qb_PM2 qs_PM2 qinv_PM2 qdef_PM2 gcrg_PM2 gtau_PM2 gmbs_PM3 gm_PM3 gds_PM3 vdsat_PM3 vth_PM3 id_PM3 ibd_PM3 ibs_PM3 gbd_PM3 gbs_PM3 isub_PM3 igidl_PM3 igisl_PM3 igs_PM3 igd_PM3 igb_PM3 igcs_PM3 vbs_PM3 vgs_PM3 vds_PM3 cgg_PM3 cgs_PM3 cgd_PM3 cbg_PM3 cbd_PM3 cbs_PM3 cdg_PM3 cdd_PM3 cds_PM3 csg_PM3 csd_PM3 css_PM3 cgb_PM3 cdb_PM3 csb_PM3 cbb_PM3 capbd_PM3 capbs_PM3 qg_PM3 qb_PM3 qs_PM3 qinv_PM3 qdef_PM3 gcrg_PM3 gtau_PM3 gmbs_PM4 gm_PM4 gds_PM4 vdsat_PM4 vth_PM4 id_PM4 ibd_PM4 ibs_PM4 gbd_PM4 gbs_PM4 isub_PM4 igidl_PM4 igisl_PM4 igs_PM4 igd_PM4 igb_PM4 igcs_PM4 vbs_PM4 vgs_PM4 vds_PM4 cgg_PM4 cgs_PM4 cgd_PM4 cbg_PM4 cbd_PM4 cbs_PM4 cdg_PM4 cdd_PM4 cds_PM4 csg_PM4 csd_PM4 css_PM4 cgb_PM4 cdb_PM4 csb_PM4 cbb_PM4 capbd_PM4 capbs_PM4 qg_PM4 qb_PM4 qs_PM4 qinv_PM4 qdef_PM4 gcrg_PM4 gtau_PM4 gmbs_PM5 gm_PM5 gds_PM5 vdsat_PM5 vth_PM5 id_PM5 ibd_PM5 ibs_PM5 gbd_PM5 gbs_PM5 isub_PM5 igidl_PM5 igisl_PM5 igs_PM5 igd_PM5 igb_PM5 igcs_PM5 vbs_PM5 vgs_PM5 vds_PM5 cgg_PM5 cgs_PM5 cgd_PM5 cbg_PM5 cbd_PM5 cbs_PM5 cdg_PM5 cdd_PM5 cds_PM5 csg_PM5 csd_PM5 css_PM5 cgb_PM5 cdb_PM5 csb_PM5 cbb_PM5 capbd_PM5 capbs_PM5 qg_PM5 qb_PM5 qs_PM5 qinv_PM5 qdef_PM5 gcrg_PM5 gtau_PM5 gmbs_PM6 gm_PM6 gds_PM6 vdsat_PM6 vth_PM6 id_PM6 ibd_PM6 ibs_PM6 gbd_PM6 gbs_PM6 isub_PM6 igidl_PM6 igisl_PM6 igs_PM6 igd_PM6 igb_PM6 igcs_PM6 vbs_PM6 vgs_PM6 vds_PM6 cgg_PM6 cgs_PM6 cgd_PM6 cbg_PM6 cbd_PM6 cbs_PM6 cdg_PM6 cdd_PM6 cds_PM6 csg_PM6 csd_PM6 css_PM6 cgb_PM6 cdb_PM6 csb_PM6 cbb_PM6 capbd_PM6 capbs_PM6 qg_PM6 qb_PM6 qs_PM6 qinv_PM6 qdef_PM6 gcrg_PM6 gtau_PM6 gmbs_PM7 gm_PM7 gds_PM7 vdsat_PM7 vth_PM7 id_PM7 ibd_PM7 ibs_PM7 gbd_PM7 gbs_PM7 isub_PM7 igidl_PM7 igisl_PM7 igs_PM7 igd_PM7 igb_PM7 igcs_PM7 vbs_PM7 vgs_PM7 vds_PM7 cgg_PM7 cgs_PM7 cgd_PM7 cbg_PM7 cbd_PM7 cbs_PM7 cdg_PM7 cdd_PM7 cds_PM7 csg_PM7 csd_PM7 css_PM7 cgb_PM7 cdb_PM7 csb_PM7 cbb_PM7 capbd_PM7 capbs_PM7 qg_PM7 qb_PM7 qs_PM7 qinv_PM7 qdef_PM7 gcrg_PM7 gtau_PM7 gmbs_PM8 gm_PM8 gds_PM8 vdsat_PM8 vth_PM8 id_PM8 ibd_PM8 ibs_PM8 gbd_PM8 gbs_PM8 isub_PM8 igidl_PM8 igisl_PM8 igs_PM8 igd_PM8 igb_PM8 igcs_PM8 vbs_PM8 vgs_PM8 vds_PM8 cgg_PM8 cgs_PM8 cgd_PM8 cbg_PM8 cbd_PM8 cbs_PM8 cdg_PM8 cdd_PM8 cds_PM8 csg_PM8 csd_PM8 css_PM8 cgb_PM8 cdb_PM8 csb_PM8 cbb_PM8 capbd_PM8 capbs_PM8 qg_PM8 qb_PM8 qs_PM8 qinv_PM8 qdef_PM8 gcrg_PM8 gtau_PM8 gmbs_PM9 gm_PM9 gds_PM9 vdsat_PM9 vth_PM9 id_PM9 ibd_PM9 ibs_PM9 gbd_PM9 gbs_PM9 isub_PM9 igidl_PM9 igisl_PM9 igs_PM9 igd_PM9 igb_PM9 igcs_PM9 vbs_PM9 vgs_PM9 vds_PM9 cgg_PM9 cgs_PM9 cgd_PM9 cbg_PM9 cbd_PM9 cbs_PM9 cdg_PM9 cdd_PM9 cds_PM9 csg_PM9 csd_PM9 css_PM9 cgb_PM9 cdb_PM9 csb_PM9 cbb_PM9 capbd_PM9 capbs_PM9 qg_PM9 qb_PM9 qs_PM9 qinv_PM9 qdef_PM9 gcrg_PM9 gtau_PM9 dc_Ib acmag_Ib acphase_Ib acreal_Ib acimag_Ib v_Ib p_Ib current_Ib capacitance_C0 cap_C0 c_C0 ic_C0 temp_C0 dtemp_C0 w_C0 l_C0 m_C0 scale_C0 i_C0 p_C0 sens_dc_C0 sens_real_C0 sens_imag_C0 sens_mag_C0 sens_ph_C0 sens_cplx_C0 capacitance_C1 cap_C1 c_C1 ic_C1 temp_C1 dtemp_C1 w_C1 l_C1 m_C1 scale_C1 i_C1 p_C1 sens_dc_C1 sens_real_C1 sens_imag_C1 sens_mag_C1 sens_ph_C1 sens_cplx_C1 capacitance_C4 cap_C4 c_C4 ic_C4 temp_C4 dtemp_C4 w_C4 l_C4 m_C4 scale_C4 i_C4 p_C4 sens_dc_C4 sens_real_C4 sens_imag_C4 sens_mag_C4 sens_ph_C4 sens_cplx_C4 capacitance_CL cap_CL c_CL ic_CL temp_CL dtemp_CL w_CL l_CL m_CL scale_CL i_CL p_CL sens_dc_CL sens_real_CL sens_imag_CL sens_mag_CL sens_ph_CL sens_cplx_CL 
