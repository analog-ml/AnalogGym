.param MOSFET_0_8_W_BIASCM_PMOS=0.813523143529892 MOSFET_0_8_L_BIASCM_PMOS=1.1884464770555496 MOSFET_0_8_M_BIASCM_PMOS=11
.param MOSFET_8_2_W_gm1_PMOS=9.732784301042557 MOSFET_8_2_L_gm1_PMOS=0.7527313977479935 MOSFET_8_2_M_gm1_PMOS=42
.param MOSFET_10_1_W_gm2_PMOS=2.174540728330612 MOSFET_10_1_L_gm2_PMOS=0.8160810619592667 MOSFET_10_1_M_gm2_PMOS=7
.param MOSFET_11_1_W_gmf2_PMOS=9.002557009458542 MOSFET_11_1_L_gmf2_PMOS=1.4720347747206688 MOSFET_11_1_M_gmf2_PMOS=101
.param MOSFET_17_7_W_BIASCM_NMOS=0.7763814926147461 MOSFET_17_7_L_BIASCM_NMOS=0.5864164680242538 MOSFET_17_7_M_BIASCM_NMOS=47
.param MOSFET_21_2_W_LOAD2_NMOS=8.522806957364082 MOSFET_21_2_L_LOAD2_NMOS=3.7058304250240326 MOSFET_21_2_M_LOAD2_NMOS=11
.param MOSFET_23_1_W_gm3_NMOS=2.80293807387352 MOSFET_23_1_L_gm3_NMOS=2.6303282575681806 MOSFET_23_1_M_gm3_NMOS=4
.param CURRENT_0_BIAS=4.407831549644472e-06
.param M_C0=4
.param M_C1=6
